&         CONCEPTL�� ��    C o n c e p t D r a w   V    C o n c e p t D r a w   V   �   �����      S e a r c h   r e s u l t s   f o r   " i d e f 3 "                    1 5 . 0 . 0 . 3 9 2 ��       �   �����          TM ����TM    gI-      E-  ����R-     O b j e c t           �?�   !   !                                                   "G]###j]G"                                                        ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�ZZZ�]]]�[[[�bbb�zzz�������������zzz�bbb�[[[�]]]�ZZZ�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�����������������������������ttt�vvv���������������������������������������������vvv�ttt���������������������������������jjj�]]]�]]]�������������������������ooo�������������������������������������������������������������ooo�����������������������������lll�]]]�]]]�����������������ggg�����������������������������������������������������������������������������ggg���������������������mmm�]]]�]]]�������������WWW�������������������������������������������������������������������������������������UUU�����������������nnn�]]]�]]]���������UUU���������������������������������������������������������������������������������������������eee�������������ooo�]]]�]]]�����xxx�����������������������������������������������������������������������������������������������������uuu���������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�\\\�ccc�������������������������������������������������������������������������������������������������������������aaa�����sss�]]]�ZZZ�������������������������������������������������������������������������������������������������������������������������uuu�]]]�^^^���������������������������������������������������������������������������������������������������������������������jjj�vvv�]]]�bbb���������������������������������������������������������������������������������������������������������������������fff�qqq�]]]���������������������������������������������������������������������������������ttt�����������������������������������������iii�]]]�������������������������������������������������{{{�������������������������������������������������������������������������ggg�]]]�����������������������������������������������������������������������������������������������������������������������������hhh�]]]�����������������������������������������������������������������������������������������������������������������������������ggg�]]]�����������������������������������������������������������������������������������������������������������������������������ggg�]]]�����������������������������������������������������������������������������������������������������������������������������hhh�]]]�������������������������������������������������������������uuu�������������������������������������������������������������iii�]]]�}}}�������������������������������������������������������������������������������������������������������������������������qqq�]]]�ZZZ���������������������������������������������������������������������������������������������������������������������]]]�|||�]]]�___���������������������������������������������������������������������������������������������������������������������vvv�����]]]�ZZZ�rrr�������������������������������������������������������������������������������������������������������������ttt���������]]]�\\\�kkk�������������������������������������������������������������������������������������������������������������rrr���������]]]�]]]�����fff�����������������������������������������������������������������������������������������������������hhh�������������]]]�]]]���������������������������������������������������������������������������������������������������������|||�����������������]]]�]]]���������xxx�����������������������������������������������������������������������������������������������������������������]]]�]]]�������������jjj�hhh������������������������������������������������������������������������������������������������������]]]�]]]���������������������qqq���������������������������������������������������������������������sss�����������������������������]]]�]]]�������������������������eee�������������������������������������������������������������fff���������������������������������]]]�]]]���������������������������������```�zzz�������������������������������������{{{�bbb�����������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�ttt�lll�ggg�ccc�YYY�WWW�^^^�WWW�YYY�ddd�jjj�sss������������������������������������������]]]�fH  ;   H  ���������  ����3  �  ��������^  ��������� t    O b j e c t *   O b j e c t [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] �  �����  pm       @o@     @o@              `��@ �����
�@    �B  J          �?    @_@�d  J          �?    @_@ iu                 @o@            @o@ j�   ���� ���� � �          ��  ����&  �  ��������p�  ��  K            S    @o@�#  K            S    @o@         �N  J          �?    @_@�p  J          �?    @_@    ��  J          �?    @_@��  J          �?    @_@ i�  ��  @   ~    �q�H7@�q�Vl@  ���T@  ���d@     q)      �      
  ��% % %                   rZ                                            O b j e c t   S t a t e   L a b e l s�      @@   @@   @@   @@ �       �B      ��                        {�                           ��        |&                                        %4  �����   �=      �Q                �f              ������     I D E F 3   o b j e c t   s y m b o l 9�  �����     O b j e c t         ��      ��         <�  �����   =  ����                        �?      �?                ?)  ����)   C^  ��������                              �?        t�           ��U U U          �?u�    ��  ��� � �         u�    ��    ��                                   m3       n)  ��  k                �!  k          �?    @_@n/  �E  j           @o@�g  j          �?    @_@��  j          �?    @_@��  j                ��  b         �?      �?        U     �?�  b         �?      �?        V-DT�!�?ݕk��|�?X���x�?n3  �L  b                  �k  b              @_@��  j          �?    @_@��  j           @o@��  b         �?      �?        U     �?�  b         �?      �?        V-DT�!�?ӕk��|�?Y���x�?&H  ��������2       �E-  �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  ^IDATx�	pTE�_��M@�(��W@!�"+� ��ˑdQ��tU��Z\)VЭB�`K֪�uK�t%���%*,��"jB���\rL&w��o�'a&3o2��W��7�u���������_wk�:����"Y�6��ѣk}}}���莜���Ʀ��ť�;1***��8W󬒿���곜�q_���w�رc'8P�uDC����4 skbb�������ڵj�ʒ��VסC��֭[ǵi�&>%%E#�f2�4�h555ᵺ�:�l6k�/_��t�R��s��Ξ=s��դ����-������~φ�F+w�}�uIII��o"_n���۷oe�޽S�v�ӭ[7�5���D�dо��[�ĉueee�Ç'@�K���b��uӦM?��eAH �H0eʔ��%?�Wއ�jذa�����:w�Q�L��C;u�V\\��ݻ�Jii)�E|)5�k�c-�4%aqNj^���x�?A�=��[o����N�߿��:�2Y�G�&�o��v��eٿ4M�!�BB�j��Ї	�,	 �3
�� �(w�T��(z!�+�(�����h��
�!�)Wq�y?�H ��P장����ѣ� ?^��p=D��U;v�h@�؈b�2�RyB�h���������7f̘��P�U���m۶�n�����[�q,�wQ֢D}9�$��o�B�<��>q��8��؄�/���������������.�f�̜�QS�N�}�?�1�4}��H��݁*5CAAA��\���5k���8����yPH@՟I��Vǎ{<��#)7�x�?�i~��w�K/�d>}��1��_�D�:�1~aԴiӞ��_y�}�uz衇��8��:)��w�G-�[�l���_���@�2`5A^^^������?���m۶d9��]/^Ԗ.]ZN��6������"��	P�r��?�4iR���>j��_�t����1��=ztf�ϰHדFH���_8c�KII	eS��y��D~��o5���֭��f/Y�$��ʟ7 �o�^9r�����Cz��93t�D�7i���P���ԩ����/N�p��܉l�
cl)?��i��m�-��`������Q�F���O�q{ux/
>|�	��+�ɩ��f(��}����)B&Lh��Ɨ�ƍ�r����c����n	���K*Dx��9_6>#�4X�.�;6�IwIU�`=�ʕ+����ddd��R�6�|B����9���͛��{U/%p�-�DcfN��i
���#G�Tz��=Z�I����g��ɓ�ϙ3'Ξ����*�P$3�����ߎ��"'ؖ~�Q� k�} r�����	3��̙i8Ŋ����|jQM@ۿ<===w��ɾp��^$ƌ9t�PL��1�?t���J�k0�Ǡv�%ɑ<��`O><��}����z�*��ѫH�H��O_���,Z�(�6)�U�p!p�n��&~	w�n_������.o�&]�8���gϞ����.E��]w�֮]�X�����
V�:=o�=3�@W�A�q�dL��'������/���R���a�|��"�T��B8��"�Nz��1	H8���,�H��z�찂��#8	^���cP�<�= =�ӴU� H@��/O_�	�1����>��j<�l�ộD�q���I6<"Ajj����x�<IS�	�d��%�y��$`L`,m� Fuw'=ɀ
�	0�/3�����nI@B�9sf�2�eh=�7l:/��Y�$�E�u2d��t�����&�	��e�Y0&��Y�f�4��z����r��g�`ZVVVs�ճ���'8
����8�>CDU��\�OWYvJ"�a�D��]�S��H���)�:˶S`mz��#��G�Ld�wOp<Wg����E���f��/�LbazO�\ߦE���w�:�,�TT��[�\!�ئ%���fegg{р�R��߂+&�YM�ӈJ`���n���������I���ӈ��;��`+xp��#D���+8;�	pF���Q1�QBv-�
Ύ�jD&>��iN��udI@��Ke��C:��VL&q|��#L���̚��%��$`9�����FX�Uq�H��*��|2���NƝs�\�l����,xۊh'k���@M&�I&��LP��g�[m$�b��]�t��W���,"����[I�R��Pc5��.�*�M4xW1���ܳ� �0v(��&%�oz	V�t[sН�f� C�%��"+	�z��"��h!x�_��N~�VC�b E�-�0�DƘ�d֊:�#�[p��öj��q %��X����u�Z��cc�@�ܥ�VP-��K
/��-��I@��=E#�B6�F$���`$��?���X�!��6^Ƒ �����gBttJ�����|	ޘ����HP+�<��8�����
\͍#URq=�w��&��e6SP�1�o��N��l�j ��
ނ��h�߫��X����������O}c�Ð��w;	�����J�!%b�B����n�F$���|�5�D����b�=�ej �4��5�{�wVT�?�@b0nQ/\���w��n'�\0�Tr��I�J�@%?q��mU
��Vc�\TTTlc�5� �Cp�mŴ���'l�f�=P�ȕ��,x�Jh'7��,$�!e�h"�,�
΂���v�]�֌r;jٞ�sJ@��o[��$�tֲ�f��:G����*�u�%kD��7}��������>��
��F�b5"Aaa���]Ŷ�a�u�H@p|g�"5"�<@qX�{�n�f�(��޳gO�4-�5$@/Xɾ��Ih*����G�PT��iQ�!�T���ꫯ��U��X�ĥ������ݴא@�n��e�{�i$�;�$����-�rg9wE��/��2��e���x�^I@p<4Z�,�NI@-p���2)gR�{7n�Ʃ� �ӯ�)	�������)̊���(���@p|���K���g�Yt�X�]oݺ��
�����l6?I�̌���!,�mݺu5�����,	�NF��ġ�G�I1D�	n����\�%�D�?}�;�S{�����Q�BL?���&�	~��$�-lziŊw���#�7�|�"�	~�r�� =�get�ȑ#��S�C@���E-�GO��	P���˗��u<k��>������z4��#H��21'�m3xETov'��G�
݅�=�����L�OG���W����"�Nz����0�f�q�ҥK˕%Q���V�\�I�c�����Ň�s0w1c�С�%������^/�����CE�W�^�7u�$��m�v3���			��TIWm�7�*�{	l޼���Ij�q|����^�k׮JV��r�JKYY��\�~��ȟ���/��ye���&�>|�R߾}��ݻ7�=xMj�l���2a�dm���j�<p�e@7�&��K�s,33�a�ȑ#����u걯$ k-X��B���o��h��w���2f��"�b��1bD�,���J }L[�h�����Z�jYK��bHpb�޳gϮ�n�{��+"��f��'�͚5KL��(((x����y4cƌW�^��5������h�7o^�ܹs�a����̸q����4���U#�ン� O?���!��^���� I{>%��J��nFF���|���C��Sn�e���,#�p��r��y�&�a�r��$��@���,;v����ejӦ��׫��$ �!���?�>�.�7��B���}�5�x�_�MOOW�q�D�9��˖-Cнk֬�����	$��S�Yy�B�K�L7�|s,�<ΜQ�O�o�Qɰ�y���c�" _'=���º�]�v�͟??�-y�Y��N[��|�f��}`2�@�F¶�S�N}t�����
u��>EBz"���)� �&p,Pnnn&�s�g����ٮ���ٳg�_|�̂Rߡ �oذ�$�2	8	~,\��iӞ`f̳&L��8q�Ɉ��� ���X����Y�_m>X$�r]!;�ːaԜ9s�pR��V��]4]ڧ�~������C�ô�'��^�?Gq|{BgLϭ�:K~/��i�	�Jo���������yAH����ɓ'O�/�����O6l�l�b{�gك��v��`W��I��t��B�@!E��~���[��?~|¨Q�b�qCoҴ?���u*�����=d���P!��#I`�O^^�-�����$�ϵ999)��P��Y=�v��i�,{P���߲����!M�|�A���p/��Chԙ���18�4`� ���,hg�w/�X(Ҳo�>�w�������Y@A�</8
�ڡ#z�d|�!��ݻw�P;���1�O�>�n�cp�\�С�����e_���Ǐ'A��|���_����/�ԑhؑ��l�*�ne��� �H�I��[�nQ�Y$c��cT�4ot
��Cιs�4��g�g9�zh�	�^���[�-�+O_���:�I�Th��ٱ �	1@�,���uw���jb�D5:F-�H=��(�!�Oc���;�>{�Gӆ���G�SC:��8�$��\�%�����o��P��?���JuH�;    IEND�B`�   g4f      0f  ����=f     I n d i v i d u a l           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�\\\�ZZZ�]]]�```�^^^�[[[�]]]�___�___�YYY�[[[�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������___�������������������������������������lll�sss�������������������������������������jjj�]]]�]]]�����������������������������lll���������������������������������������������������������kkk�����������������������������lll�]]]�]]]���������������������bbb���������������������������������������������������������������������lll�������������������������mmm�]]]�]]]�����������������jjj�����������������������������������������������������������������������������rrr�ooo�����������������nnn�]]]�]]]�������������UUU�����������������������������������������������������������������������������������������|||�������������ooo�]]]�]]]���������fff�������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�����eee�����������������������������������������������������������������������������������������������������kkk���������rrr�]]]�]]]�����������������������������������������������������������������������������������������������������������������ggg�����sss�]]]�\\\�___���������������������������������������������������������������������������������������������������������������������uuu�]]]�ZZZ���������������������������������������������������������������������������������������������������������������������kkk�vvv�]]]�]]]���������������������������������������������������������������������������������������������������������������������iii�ppp�]]]�\\\�������������������������������������������������������������������������������������������������������������������������ggg�]]]�����������������������������������������������������������������������������������������������������������������������������ggg�]]]�����������������������������������������������������������������������������������������������������������������������������ccc�]]]�����������������������������������������������������������������������������������������������������������������������������___�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������aaa�]]]�����������������������������������������������������������������������������������������������������������������������������fff�]]]�vvv�������������������������������������������������������������������������������������������������������������������������iii�]]]�XXX�������������������������������������������������������������������������������������������������������������������������ppp�]]]�___���������������������������������������������������������������������������������������������������������������������]]]�|||�]]]�ZZZ���������������������������������������������������������������������������������������������������������������������uuu�����]]]�\\\�ccc�������������������������������������������������������������������������������������������������������������lll���������]]]�]]]�����ttt���������������������������������������������������������������������������������������������������������������������]]]�]]]�����vvv�����������������������������������������������������������������������������������������������������ccc�������������]]]�]]]���������ddd���������������������������������������������UUU�kkk�����������������������������������������UUU�����������������]]]�]]]�������������UUU�������������������������������������UUU�UUU�UUU�������������������������������������]]]���������������������]]]�]]]�����������������eee���������������������������������UUU�UUU�UUU�xxx�����������������������������ggg�������������������������]]]�]]]���������������������|||�vvv�������������������������iii�UUU�XXX�����������������������������fff�����������������������������]]]�]]]�����������������������������bbb�����������������������������������������������������^^^�������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�rrr�iii�eee�YYY�xxx�������������������������]]]�aaa�kkk�}}}�������������������������������������]]]�f Q  5    Q  ���������C  �����C  � x 
   I n d i v i d u a l .   I n d i v i d u a l [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] �?  ����	@  p�?        @o@     @o@          �������@ VUUUUu@    ��?  J          �?     @_@��?  J          �?    @_@ i�?     0���2��     @o@"+?!�Mh�    @o@ j�?   ���� ���� � �          �B  ����sB  JA  ��������pA  �J@  K            S     @o@�t@  K            S    @o@         ��@  J          �?     @_@��@  J          �?    @_@    ��@  J          �?     @_@�	A  J          �?    @_@ i(A  �&A  @   ~   �q���E@��8���i@  ���T@  ���d@     qzA      �      
  ��% % %                   r�A                                            I n d i v i d u a l   L a b e l s�A      @@   @@   @@   @@ �       �B      �B                        {BB                           �BB        |sB                                        %�B  �����B   ��B      ��B                ��B              ������B     I D E F 3   i n d i v i d u a l   s y m b o l 9-C  ����-C     I n d i v i d u a l         � C      �-C         <;C  ����;C   =xC  ����xC                        �?      �?                ?�C  �����C   C�C  ��������                              �?        Q  ��������Q  ����Q     f�K  ;   �K  �����K  1I  �����K  I  ���������H  ���������            _E  ����mE  pE  �GD  C        @o@�sD  K	            S    @o@         ��D  J          �?     @_@��D  J          �?    @_@    ��D  J          �?    @_@�
E  J          �?    @_@ i*E  �(E  A   ~               @o@            @o@ j_E   ���� ���� � �          �GG  �����G  �F  ��������pvF  ��E  K            S    @o@��E  K            S    @o@         �F  J          �?    @_@�%F  J          �?    @_@    �KF  J          �?    @_@�mF  J          �?    @_@ i�F  ��F  @   ~       @_@    @_@  XU�Y@  TUEb@     q�F       �      
  ��% % %                   rG                                              s@G      @@   @@   @@   @@ �       �B      �GG                        {�G                            ��G        |�G                                        %�G  ���� H   ��G      ��G                ��G              ����� H      9/H  ����/H              �"H      �/H         <=H  ����=H   =zH  ����zH                        �?      �?                ?�H  �����H   C�H  ��������                              �?        t�H           ��U U U          �?u�H    ��  ��� � �         uI    ��    ��                                   m�K       n�I  �^I  k                ��I  k          �?    @_@n�J  ��I  j           @o@��I  j          �?    @_@��I  j          �?    @_@�J  j                �>J  b         �?      �?        U      �?�vJ  b         �?      �?        V�!3|�@ݕk��|�?X���x�?n�K  ��J  b                  ��J  b              @_@��J  j          �?    @_@�
K  j           @o@�BK  b         �?      �?        U      �?�zK  b         �?      �?        V        ӕk��|�?Y���x�?&�K  ��������2       fQ  ;   Q  ��������IO  �����P  1O  ���������N  ��������� q         �L  ����zM  p�L  �L  G         �A@      �A@         �JL  N          �?     @_@�rL  F     �������?    �m@    ��L  J          �?     �1@��L  J            �A@ i�L                  �A@             �A@ j�L   ���� ���� � �          �                     {IM                            �IM        |zM                                         %�M  �����M   ��M      ��M                ��M              ������M      9�M  �����M              ��M      ��M         < N  ���� N   ==N  ����=N                        �?      �?                ?KN  ����KN   C�N  ��������                              �?        t�N  ��N  F                ��U U U          �?uO    �� ��N  F      - ��U U U ��N  F           �O  F        u1O    ��    ��  �)O  F                                       m�P       n�O  �vO  k                ��O  k          �?     �1@nHP  ��O  j            �A@��O  j          �?     �1@� P  j          �?     �1@�P  j                       �?         f�k��|�?T���x�?n�P  �eP  b                  ��P  b               �1@��P  j          �?     �1@��P  j            �A@       �?         u�k��|�?G���x�?&Q  ��������2       Q  ��������    q � Q    �0f    �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  qIDATx�p�ն�w:�H�Q0��!��irA@Ј�}��R��#2�SG�Q�\�>y
H���t��J�&҉`("�	!y�u�䞄S�ӒsN��9�����o��Z{J�_��@P s`���!!!����	

�\�5�s?���8�c>������/��2��p~255�<��:�yIII�jժ%���u,((H�:�F��u��-�馛�8��^�zhDD�
U�S D���"����/�_���Ux����K�.E\�vM��=���� �n��^�dI^  �oA��C5�M���>::�z˖-�n�������n�M���y��$gϞU�O�V�N�*8x�`��s�"##�Q�J@�5}(�{��
.į@0x��v0~8��(oblbb����5k�x�+�u��Ǐ��{��ڵ+'##��&|-�bNnn�j~� 7*�y ����Gt?����޽{D�.]�n��7��|V��c��aÆ�H�p��T���<_�gK�Y2�"~�����[ܷo��ƍ{�z/�����֯_}�ʕ�H�H��rrr���t�51���'��߂�����9�Rwy�X��lٲ��G�����w�ʕ�!��5��g@@����׮];>%%�4ޣ����S�����˗�n߾�0��l�}��l_hv�sY�=4��������Ǣ��_��fj��9���+Dgxa�ҥ���\i 4hP�����s�O<ѳg�`�m�d'O�T3g�̾p�Bz^^��*S��<��Ï����ݻw8�՘�DǺBĶm���ٳ�"�"^��!�BAп��X�aĹ�g��NHHp�o�ۂ�3gN��ݻ��I�L��"��0���Ř��_�~��<�H��k��,��{ｗ{���(��lܸ��l
�\U�{챷���}��[�h�J�T��>��y���+Vdx�4�����&s��4h7q��hfަ'`�_�xq! ��ؔ���ݛ�yM&3�o v��5}��g#�s��9�3,�Q�F�iii)M�6=q�С�s;��+ @t�ӷ0��� ,��>α׽����S:t��ԯy��a?���&�J���� ���	���?VL�֫�w�r@���0c搈D�����F�M�Q�@ ��ŤI���4ib�:�`PR�F�*>{�ܹO�b8���T������(� ��o<��f͚��m����=jj��p����v̘1a�۷7N�N� �B�!��	��������>k�۵k�Q:�� t��5|�֭-	����� @�Զ�c�Ƶi�ƣ����:9$H�cǎ�D1u nO]A�>}���������\N��:�R*:CoئM����܀!��\V	�^��~rrr����|�q�~���瞋�'��5���<lذ�D =9ah�r����'%��B��d�C�k��%;Q�	̛2eJ4A!�֧�{�bbFA�b�1�u�
������=ztd�Z���K��"ƍ'Ry,/��V����VZ�S�Nz&�,������@^�TwN�k�@�RF��ezt�.r�i��Ȋa���L�@����a�9S�N[�����ߐ�Vmh�/T���ru�J���h9�h�@��\���/G�8�h�:]%r@�i�\��o�#�^GMq(	@�t�CC�ԩ�,�܇8��SO�n0͈�h,iʆ9��}�)8@h�BQ����8Jn��2+�ʠ#6��s,��(�P����a��A��o�7;�H��	6�`���	����a8'����|��)�s2ͷ�T� @��z(�le������P��R��b�  \|�%�Ad�m�u��=�n��V[A��<�@�]*l�[~z/�bX�cˊx퍇0\��8@��lPm�5�n c�h2�@k���{=z�A�lMA,I��$|�U��n�鲒�>���?/��
+zc������ �����K/P�ҭ[7�֥��k���=��#�8�BA,�8�AcF߶m��U��Nq@�����d��2c)�܅���BK��9�^4���jIY)��Nh��Zr' ϑ��m�%i� @
$�q����%U��&X��X枀^Pj,
CG@`3�~� �E�!�t�X|��['��Z���hGT`F�O�� h���B��s�@����h����\�I���lz�c��\	�㭷ު�F�.3�&�/H�R�gf��Q���vS3�f�0�U��{�����P=!�>1�@���ˑ�K_�`�;2 �Ӓ����}�S�P��_P� �d��B���rh�_@��Z(�ת��T8�R���?@@8rMP�_�Խ�: �|e��D�)�H"���9e<$�i3d��_��:���ah������/s���� `8(a�_��:�"JfS���%��s�#�s�˟/m��Pm&�ǎt��؇��B�w��y����H�ߤ��r��˄ �!M��Nr��իE� ���c#��W9�&N2�ߓ_�r� ��%�#�o�]E������w�|xS\%�(��l�ү��*��WE8@��rM `��i>�^E��d
� �	97���������Tb�3�YB�	(�i'N�ȭ,�T�a�*�cfN�@ *�;vL�����3g�(,�;�d�@��`?�B$S�}}`?~<;???�L�	�W��d��!bB��,A�o3Sj�\ 6���O�����R�rrrB�6�X
�=p�@���>&�EG)�7ԕ��� @�ٷo_8����^Se���ݻs��Y������	9:���?[>��Ɓ��4���$�r�i�{���NK�9�T:�lٲ2oz0mX�~�zS�I ѮI��[�l��XX�!e@ B���$WO˳)0�7n�X@��/OM�C��<����s�ϯq($}6���I�������:��<�����o�ɣogZ��`D8�k��h��@��[�#��e��@ �����]�r�6Y������	#��n5r�*._����ɓE���d�dK�S����"<���U�E1~���c�X��dXg88�t��-�Zo����ܳgO��=��:���hѢ,��${��		=°0u��:��}�~u�ҥ�?���i��i��~���_~�W�~����OE
ȇ1K=�֚j(� �>��lk��=����u�Y[p)�V��d������+HGe��>�L�j޼y����H��@f
:J���"ai�Y�x�8�[3[k�CH&��������ָ�C��W��1��5�,C ��(���~�m��0emŧ�,����l<�����F[`z��̣�}��l*1Z�NW�����X]������{�0)���*Y��'���{\��g�R�V��c�a���;)�a�6oޜ�gβ�{��iӦ� ��ꫯL{8S�K[��)�D>����ߎ�{:��W�ie1�;����Ś&6�5j�&M�(�x$_��6:� ��WrXZ6��>{ٙ��.�@2����dg�i�1ı���٣(ML��p����v�Y@��O*��}�ܹ�v͟?�Dٵ�":��G�Y���f͚%plڵk�p�Hu��Ҟ��Z���;
�����mǹs��u�E��f͚v�V��5k�\_�|y��N��j{\�TV2�ªX�7�'��q9}�t���<I�k�.թS'����UdB<�j֬YYx{;a�9�N�n� ��0��2��1q�Z��9 `8QDI9�#�d	7w:��3�L`�ԩ�>  ~t�>�@ ������#ңXc ��e�K�9��~�%��[Ne���͛+_�4� ��^o? ��)�l$��@���7<V��Ǝ�3��a����no�V���X/��Ť� X穪<i��O/^����Ӿ�c8|�t�����D.Wn���ѣ��7��%f�����>��%h�H��D6�81s��|G��ۭwP�o��vmu���c,p�T�ӝ;w�L�<YvIF��t��4N��AG2;�x�{srOS�<OL[�ѣ|�z�R[4cƌ+Ls���ި�� �FJ|"��E0���Ǐϖ�we�<1ϯ��������)t
����� W��5M^���fW4n���z�}�0���J]�#���]�/;w����n�e43�>ԫ����S����������a��k 0W"�E��k�q!�[�e����W�"	pv�=.�3bĈ
�n߾�dʔ)y8�^#Pt@�߾Bz��Y��
�&�p>��r��(�y\\�B�2��L:�#��߿�=o]�i{��ٹL�/�>�,�V]�˭H�G��gxX� ���v�l�2��[y�,�6l(�����Ӗ���饗^R|;�aZw�����_�MOO_�R���/�<�n����wРAu� �"##{�92�]�vδ��	��*�����x5a�U�~}��r&�X$?����'��SP��:��Si+��2$	 �nԨQ����v�Z���iE�ԫW/q����s3=~я�/`�'�շ�ELŶbۿ���-�RA M�޽{(o����:!tذaQu��-�J^�ԋ͹J�JDJHPIBB��С�W�@�[����� �r�~�cW��\܃$;,��A`n�СCc ��0�E�dA��FB���M_�_#�fߵ\�������3 03d���(cc�T�%@�������䳮������#H%��/A~�eaG|����A2L`��9D�޽{�t��%��c e�`���~v�B\���t�O	�7��kG��%�*��02=�"գG�jm۶��PoO1-�a�\�|�36mڔ��φ��y�ga���<.��٪�����K�3�E
��[vs�6m
���8[�H��p��Y����� ��+A��ֿ��U���[���߁��0��ztz� {q����"M?�T�D�_f���.o�yï��O:��(�y�w���6���]>��[���ܯA`I��'%%�1�o�ޚu���[Gm��b������Ӊ
i$�	�Kd�5�[���(�^8�3��S�1����4���-_�?_�uzEu:P�PpĒ6�D�������H��H�����ǧ�0~�~u�E�
��    IEND�B`�   g^�      Z�  ����g�  (   W e a k   T r a n s i t i o n   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������|||�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�~  <   <~  ����<~  $~  ���������}  ��������� �    W e a k   T r a n s i t i o n   L i n k 8   W e a k   T r a n s i t i o n   L i n k [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] �y  �����y  p�y  ��x  K    
   Sª���&w@         ��x  K    n���!	@   
 <        �y  B   
     %   _UUUU�y@�/y  B        %        ��@    �Uy  J          �?ª���&g@�wy  J          �?         �����l@      ��@ `UUUU��@      ��@i�y           �ª���6w@      �      @j�y   ���� ���� � �          ��{  ����r|  9{  ��������p{  �#z  E   *   �ª���&w@�Dz  M   *    X     �I@�yz  H    �'DT�!�? �'DT�!�? g        ��z  H     Zª���&g@��z  H     [      �9�    ��z  H          �?ª���&g@��z  I          �?     �9@ i{  �{  @   ~   ª���&g@ª���&g@      $@     �D@     qi{       �        ��% % %                   r�{                                              s�{       A    A    A    A �       �B      ��{       �|  ��{  H          �?ª���&g@                         {A|                            �A|        |r|                                        %�|  �����|   ��|      ��|                ��|              ������|     w e a k   t r a n s i t i o n   l i n k 9:}  ����:}  (   W e a k   T r a n s i t i o n   L i n k         �-}      �:}         <H}  ����H}   =�}  �����}                        �?      �?                ?�}  �����}   C�}  ��������                              �?        t�}           ��U U U          �?u
~    ��  ��� � �         u$~    ��    ��                                :�~  ��������                                                        �Z�  �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  :IDATx��1    �Om�@a��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`�<0� ���b    IEND�B`�   g��      ��  ������  ,   S t r o n g   T r a n s i t i o n   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������|||�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f��  <   z�  ����z�  b�  ���������  ��������� �    S t r o n g   T r a n s i t i o n   L i n k :   S t r o n g   T r a n s i t i o n   L i n k [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] �  ����%�  pړ  �В  K    
   S�����&w@         ��  K    n���!	@   
 <        �:�  B   
     %   `UUUU�y@�e�  B        %        �@    ���  J          �?�����&g@���  J          �?               l@      �@ `UUUU��@      �@i�           ������6w@      �      @j�   ���� ���� � �          ��  ������  o�  ��������p7�  �Y�  E   *   ������&w@�z�  M   *    X     �I@���  H    �'DT�!�? �'DT�!�? g        �Ȕ  H     Z�����&g@��  H     [      �9�    ��  H          �?�����&g@�.�  I          �?     �9@ iM�  �K�  @   ~   �����&g@�����&g@      $@     �D@     q��       �        ��% % %                   rЕ                                              s�       A    A    A    A �       �B      ��       �<�  �+�  H          �?�����&g@                         {w�                            �w�        |��                                        %��  �����   ���      �Ӗ                ��              ������     s t r o n g   t r a n s i t i o n   l i n k 9x�  ����x�  ,   S t r o n g   T r a n s i t i o n   L i n k         �k�      �x�         <��  ������   =×  ����×                        �?      �?                ?ї  ����ї   C�  ��������                              �?        t*�           ��U U U          �?uH�    ��  ��� � �         ub�    ��    ��                &                :��  ��������                                                        ���  �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  :IDATx��1    �Om�@a��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`�<0� ���b    IEND�B`�   g��      ��  ������  4   n - P l a c e   1 s t - o r d e r   R e l a t i o n           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�[[[�UUU�}}}�������������������������������������UUU�___�\\\�UUU�������������������������������������������������������������������������������������������������������������������������aaa�YYY�YYY�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������ZZZ�XXX�����������������������������������������������������������������������������������������������������������������������������YYY�]]]�fff���������������������������������������������������������������������������������������������������������������������UUU�[[[�\\\�bbb�^^^�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�ddd�eee�eee�eee�fff�jjj�ttt�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�fO�  ;   O�  ��������e�  ����:�  M�  ���������  ��������@�     n - P l a c e   1 s t - o r d e r   R e l a t i o n >   n - P l a c e   1 s t - o r d e r   R e l a t i o n [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] ȭ  ����֭  p��   ������r@      @_@          �M6�@ ΡbA�˕@    �`�  J          �?������b@���  J          �?     @O@ i��             ������r@             @_@ jȭ   ���� ���� � �          ���  �����  	�  ��������p߮  ��  K            S������r@�A�  K            S     @_@         �l�  J          �?������b@���  J          �?     @O@    ���  J          �?������b@�֮  J          �?     @O@ i�     LUUUCD@TUU՟7p@   ���D@   ���T@     q9�      �      
  ��% % %                   rj�                                            R e l a t i o n   L a b e l s��      @@   @@   @@   @@ �       �B      ���               d�  ��  C         4@ |       4@��  C   J    ��?�߾�?;�O��n@        {N�                          �N�        |�                                       %��  ���� �   ���      ���                ���              ����� �     n - p l a c e   f i r s t - o r d e r   r e l a t i o n 9c�  ����c�  4   n - P l a c e   1 s t - o r d e r   R e l a t i o n         �V�      �c�         <q�  ����q�   =��  ������                        �?      �?                ?��  ������   C�  ��������                              �?        t�           ��U U U          �?u3�    ��  ��� � �         uM�    ��    ��                                   m:�    	   n��  ���  c   J          4@���  k            @_@nV�  �Ѳ  j                ��  b    J         @Z@��  b   K    ;�O��n@�,�  b    K    +��]@       �?          ��z��?��[�V��?n��  �r�  j                ���  b   J          4@n,�  ���  b   J          4@�̳  j                ��  b   K    ;�O��n@��  b   K    ;�O��n@       �?         ML�Nz?iUVD��?np�  �J�  b    J    �����q@�h�  j                n�  ���  j       ������r@���  b   J          4@�Ǵ  b    K    ��ʡEbr@��  b   K    ;�O��n@       �?         ��Px^U�?�N)Sj�?nP�  �(�  j       ������r@�H�  b    J         @Z@n��  �n�  b    J    �����q@���  j            @_@���  b    K    ��ʡEbr@�̵  b    K    +��]@       �?         g�b��?S�=u���?n:�  ��  b                4@�2�  b               @_@&O�  ��������2       ���  0  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx��OHa��wg�/�EE�(�Y*&�Bԫ�Q�y-<t<�t<Q�B�"� "K

�J�@C�U�]��y7G��Q�����ٝ�y>�c�w���R�@ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ �����Q]]�������-�\��0<<�=J^�W�ASSS��r=�B-�X����Q����e��ﮟ@"���nw�������\__�411=��B������x>VTTx���ҋ��Uzz��߱~Cvvv�������ܖ�y=��×ӻ&�����𺣣#XPPpz;� ����:;;U x���?h�t����	�@OO���Ȱ���akkk����`oo�adddL���d�%��o�������/�
������R�����������1K�*3���՞��\��NY�
Uee�7����4���OoȲ�jkk�$�u����%�������]5՝())Q�h�Lܖ�ȖK�׎g~����6��y��������|p�%�	PPJ@�{"�RsL� f�T�����D��l�f�T���0�����@�-�p`��OUOs2���� �1 d�3`8 Z�99 d�3`8 Z�99 d�3`8 Z�99 d�3`8 Z�99 d�3`8 Z�99 d��L }�iWcf�Ҿ�e%��u�KsC�D���쏵���!M�ݲb ��%omm)�}tttߚ���K��ə�sE�|zz:)��to�d��@z��H|9�+Y�֩���}y���ۗ�_%?%1�H̫���Kr�s���S]Υ~2//���dn�)++��a���+��닇�a�������Ó腥��=i}�N�h��<��'-oNbNy�9����2�uxxX466�kW����������.�x����(//dff��^��	�7D@���܌���E766����[�e83�_�]�~�����ߗ��<	��m��.0�H��2៑I�������uv@ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ ���_�L"0��T    IEND�B`�   g��      ��  ������  4   2 - P l a c e   2 n d - o r d e r   R e l a t i o n           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�YYY�������������������������������������������������������������������������������������������������������������������������|||�]]]�UUU�UUU�ZZZ�^^^�___�___�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�\\\�WWW�YYY�XXX�������������������������������������������������������������������������������������������������������������������������zzz�\\\�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f��  5   ��  ��������O�  ����O�  � �    2 - P l a c e   2 n d - o r d e r   R e l a t i o n >   2 - P l a c e   2 n d - o r d e r   R e l a t i o n [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] P�  ����^�  p�  �	�  K    
   S��8��"w@         �H�  K    n���!	@   
 <        �s�  B   
     %       ���@���  B        %      @=�@    ���  J          �?��8��"g@���  J          �?         �qGt�@    @=�@ r�q܂�@    @=�@i�             ��8��"w@   ���F�        jP�   ���� ���� � �          �k�  ������  ��  ��������p~�  ���  C   *   WVUUUl@���  C   *    X   ��*H@���  J    �'DT�!�? �'DT�!�? g        �
�  J          �?��8��"g@�-�  B          �?   ��*8�    �S�  J          �?VUUU\@�u�  J          �?   ��*8@ i��  ���  @   ~         @VUUU�k@      @   ���F@     q��      �      
  ��% % %                   r�                                            R e l a t i o n   L a b e l sd�      @@   @@   @@   @@ �       �B      �k�                        {��                           ���        |��                                        %��  ����^�   ���      ��                ��              �����^�     2 - p l a c e   s e c o n d - o r d e r   r e l a t i o n 9��  ������  4   2 - P l a c e   2 n d - o r d e r   R e l a t i o n         ���      ���         <��  ������   =�  �����                        �?      �?                ?�  �����   CO�  ��������                              �?        ��  ����������  ������     f��  ;   ��  ������   �  ������  ��  ����������  ���������            �  ������  p��  ���  K	            S��8��"w@��  K	            S                 �H�  J          �?��8��"g@�k�  J          �?            ���  J          �?��8��"g@���  J          �?         i��  ���  @   ~           ��8��"w@                 j�   ���� ���� � �          �                     {U�                            �U�        |��                                        %��  ������   ���      ���                ���              �������      9��  ������              ���      ���         <�  �����   =I�  ����I�                        �?      �?                ?W�  ����W�   C��  ��������                              �?        t��           ��U U U          �?u��    ��  ��U U U         u��    ��    ��          ���  F           ��  F                           m��        nw�  �M�  j                �o�  j          �?        n��  ���  j       ��8��"w@���  j          �?        &��  ��������2       f��  ;   ��  ����������  ������  x�  ����������  ��������� L         J�  ������  p�  �O�  C         >@ |       >@�u�  C         >@ |       >@         ���  N                ���  N          �?            ���  J                ��  J          �?      .@ i�                   >@              >@ jJ�   ���� ���� � �          �                     {��                            ���        |��                                        %��  �����   ���      ���                ��              ������      9@�  ����@�              �3�      �@�         <N�  ����N�   =��  ������                        �?      �?                ?��  ������   C��  ��������                              �?        t�  ���  F                ��U U U          �?uN�    �� ��  F   - ��U U U �6�  F           �M�  F        ux�    ��    ��  �p�  F                                        m��       n��  ���  k                ���  k                n%�  ���  j                ��  j             >@nk�  �A�  j             >@�c�  j          �?      .@n��  ���  b                  ���  b                  &��  ��������2       ��  ��������    L ���    ���  �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  "IDATx�ֽJ�P�:���5�t�z���͸�x���p��������%�d;�	N9?��{�< @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� �����ju4�N�6�M5�Uv�*І`�X����(���d� ��sع������x|�e�I��g�03�]�!� �6��>�T�9���BнF:����eY�Eїۮ[��g�?E{޶�\z�͑# ��-��}�O nc�&�{�c�
�!���1>�n��W���z�ҷ�X�mz��?��g߆��@����;ܧ�&x�����w@��  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� :�oK�L�"�;:    IEND�B`�   g-     ) ����6 *   A N D   J u n c t i o n   ( o b j e c t )           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�\\\�[[[�YYY�YYY�XXX�YYY�ZZZ�[[[�\\\�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�����������������������������������������]]]�zzz���������������������vvv�___���������������������������������������������jjj�]]]�]]]�����������������������������kkk�������������������������������������������������xxx�rrr���������������������������������lll�]]]�]]]�������������������������ttt�������������������������������������������������������������lll�����������������������������mmm�]]]�]]]�����������������ggg�����������������������������������������������������������������������������lll���������������������nnn�]]]�]]]�������������UUU�������������������������������������������������������������������������������������aaa�����������������ooo�]]]�]]]���������hhh���������������������������������������������������������������������������������������������sss�������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�����lll�����������������������������������������������������������������������������������������������������bbb���������sss�]]]�]]]�uuu���������������������������������������������������������������������������������������������������������������������uuu�]]]�[[[�rrr�������������������������������������������������������������������������������������������������������������```�����vvv�]]]�]]]�����������������������������������������FFF�111�111�111�@@@�������������������������������������������������������������www�]]]�]]]�������������������������������������EEE�111�������������111�BBB�����������������������������������������������������ttt�www�]]]�\\\�������������������������������������111�BBB�������������444�111�����������������������������������������������������ZZZ�xxx�]]]�qqq�������������������������������������111�BBB�������������333�555�����������������������������������������������������ccc�vvv�]]]�}}}�������������������������������������KKK�111�|||���������111���������������������������������������������������������mmm�ttt�]]]���������������������������������������������EEE�111�666�333�������������iii���������������������������������������������sss�ttt�]]]�zzz�����������������������������������������===�111�111�AAA�������������111�ddd�����������������������������������������kkk�www�]]]�eee�������������������������������������555�JJJ�����aaa�111�HHH���������111�yyy�����������������������������������������XXX�|||�]]]�XXX���������������������������������mmm�111�������������^^^�111�KKK�����111���������������������������������������������ddd�~~~�]]]�```���������������������������������BBB�111�����������������[[[�111�111�111���������������������������������������������~~~�����]]]�ZZZ���������������������������������AAA�111���������������������WWW�111�999�����������������������������������������{{{���������]]]�\\\�^^^�����������������������������ggg�111�JJJ�����������������___�111�111�RRR�������������������������������������fff���������]]]�]]]�������������������������������������333�111�III���������III�888�����QQQ�111�VVV���������������������������������������������]]]�]]]�����bbb���������������������������������JJJ�111�111�111�RRR�������������LLL�111�ZZZ�������������������������mmm�������������]]]�]]]���������kkk���������������������������������������������������������������������������������������������ddd�����������������]]]�]]]�������������www�������������������������������������������������������������������������������������UUU���������������������]]]�]]]�����������������ZZZ�����������������������������������������������������������������������������ggg�������������������������]]]�]]]���������������������fff���������������������������������������������������������������������bbb�����������������������������]]]�]]]�������������������������kkk���������������������������������������������������������~~~�www���������������������������������]]]�]]]���������������������������������ddd�qqq�������������������������������������iii�nnn�����������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�ttt�nnn�ggg�eee�]]]�UUU�YYY�VVV�^^^�fff�kkk�www���������������������������������������������]]]�f��  ;   ��  ����������  ����o�  ��  ��������V�  ��������� �    A N D   J u n c t i o n   ( o b j e c t ) 9   A N D   J u n c t i o n   ( o b j e c t ) [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] ��  ������  pw�   �����V@ �����V@          VUUUe/�@ �����p�@    �L�  J          �?�����F@�n�  J          �?�����F@ i�             �����V@        �����V@ j��   ���� ���� � �          ���  �����  �  ��������p��  ��  K            S�����V@�-�  K            S�����V@         �X�  J          �?�����F@�z�  J          �?�����F@    ���  J          �?�����F@���  J          �?�����F@ i��  ���  @   ~   ������9@QUUUP@�����'@������S@     q3�      �        ��% % %                   rd�                                            & s��      @@   @@   @@   @@ �       �B      ���                        {��                           ���        |�                                        %�  ����o�   �%�      �9�                �N�              �����o�     A N D   j u n c t i o n 9��  ������  *   A N D   J u n c t i o n   ( o b j e c t )         ���      ���         <��  ������   =�  �����                        �?      �?                ?!�  ����!�   CV�  ��������                              �?        tz�           ��U U U          �?u��    ��  ��� � �         u��    ��    ��                                   mo�       n!�  ���  k                ��  k          �?�����F@n��  �=�  j       �����V@�_�  j          �?�����F@���  j          �?�����F@���  j                       �?         ݕk��|�?X���x�?no�  ���  b                  ��  b          �����F@�'�  j          �?�����F@�E�  j       �����V@       �?         ӕk��|�?Y���x�?&��  ��������2       �) �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  IDATx�	pT՚�og_	KHPdw��AA�d+�,"!�Q,�Z�+��8<3�Z�ʱ�y8�<�}��A�&P�";�E���2��!y�;ݝ�s�snխ�}��|�w��;���w��4u(	(	(	(	(	4z	�ƍ�إ`
F�3�Ehhh
���)22���dj]UUռ��"���2������
��y��"}!��s^�u�V~ii�)�9�����^�fMe��,�A _2����?66�	*.�J�nݺui۶m����$S�fʹ����'�4*��)���}޸qC+**�n޼�]�zUN��˗KϞ=³h��h'���2�������ѣۄ��=E��///�ժU�򔔔�nݺEt��IKLL�I���f�کS���9R��w߉6) t��c�/���3//��'��0Ӏ*>	U=)&&f_m�Gy�ꡇ�IMMո�C9��>|�r���Eh�����d�ڵkw�f�㷍��� 0edd��/�%��A}����߿_}�*7����k׮i_|�EՎ;�


J�y	��6\5�ִÇ����=_�|��#G�S�&�ck��???_۶m[)B�vX���g�p҈
b�!�?�R��ܹshzzz����oD�9M�����999f�<�Ƙ<�t~Hh��~��)�P�QS�L�k׮���_�Z��[�V�[��Lw3��Ƌ�6m��?
��� ;vl_���lٲͳ�>w��ڧ6����i�h*�{tE�ڲeKIC��` xꩧ����3�M�;`����������_��˗��7E4����w"��  �����=u��h���/�dɒ����ׯ�a��ͅ�&ʯ ���ƅ��g^y啘.]���_C�'MDvvv��ݻ������p�t��ߏs�����c��.m�rh5_ḹc��w�r�����"�/� �������3��/���m�Ÿ��q����n���k�g�yf^\\�{|��={���|-4_�/�ѐ!C"�>��x�=���'O����2}�A��a�����Y�-�U���j�a�=���axH��tl��'N���|���	����V?O���[u�.�@vBԡC�&r} @�s=����z �y7=�D����ڂ$��p9{U���_v���Ι3'J��ʯyo�ֵkWm׮]������g��� u�?|����
 ި��At�&C�U��w�}� ��<���[�� �6,u�ҥ�
 �U���Ź����0Ж�kO{�\��M0iҤEX����&��P��$ �s��9��<v3{\�S�4i� +++6��>|WM����{�1�q������￿�I�� O`���|��X_wz�\0�K�;����1���)����W�A�h ̞=;{��]MO�j,��߳gO["��k8�.�n������Lx��G ܕ����$ho��F,s(��V~����Z`!'O��n��=�H@|3g�d�6f�:�3\n蚴�؜��״iS�p�r�H�c����������˚�����؀�e��>� ��1�,N�Yx��b\A�h����V2ϒ@�(�V�\�����Q�b� �P����B�ͽo߾�6m�$c(>�JN� ��tI"韺��J�g	̚5+d1k���E;��尿y�������,G�<������0���YQ8�@�СCCe��:�/l�h��M�'�T4o� �� �p2*�����6��u���C03�!�^`u�e�8m�L~*�A$ -�gLB+���$� HKKkJFSG���w�O�F{.m�~�L�XmA�g���Rݼy���Q�(�9����:"�E/��P=G4�3�r�:t�`�˛�L� �;8��@�,���������ҟq`��O>�&8�^ <�ݻ�Pٕ1���ȵ	�d���
�|n/3u�x?~�дO�G��JnѢ�Ȏ;�U�О��>���ۣ�&0$�5���`�	��[�kl� ��`�>`�*rI��?YJo��4u@���7��J��%����,����lqP,�;DnŪ�*@�3�D���ro��:��ꀀ���lQnbcԝר�^54����T�L�A`b�Lx�N���X6���~֬X� _sz�kh-���ϴ�hF��Xsc��byvkF���%@��$��� F�,�Wv*E J��������$��[���e�����u`K��\�������Ģ�	#� Ӛ���~�ஃ�C�K�]
z��5��H�Y{=g�  -M�zz��5����l��D-��6�9��V�% kJ2����^-���(>�Cu|M�D�Vz�jA@;�G�����2q��"r�8�"�>Q��a��YB�ˎ��� �A$�H�Ă�]���,���jT ׳$����n�'P6�^bAx-[���[t j��5����n	H��/kA��r�KQA,�A�2=�� ��uV�T6�^:AxM�MP�g���W��ui�#}F�:0$  �'tUOm-JJJ�Zfa5����� kj����Ԃ@�^�I0�sud�r�J 8�g�r��JW�^�����:$p���rl�szV,@���,2꟫� ��|��g�lY� ���.�n�^BAt-�C6܌�C?�g�x����/�'P��#�K�.I�5//϶�@X��8�j��u<�n�ɏ?��1�x��&,楡*N0�)=������ �f���i͕Es�������u:�?$p�ر2E{�Y� �<dr��ӧO��$kI��=����Y��5+u@�#a����qh-� �ώ(��Gq
�[�ba��~�a��7o��T������W_}U�=��u4�oэ�+�QG�H�СC�6�G�a���l�D��_6'젪a�\�n�q[����F�j0ɖ��޾}�$j,��6A #��Rه
����@ؽ{��^���l�#�/[�l�i�Eu?0$p�����6l8f�b� `�)租~�W�:Wh�"��{�8��5k�T2��ann��`����3cI��������CX��G���������;wJ��(�̠ؼy�����:��9��
�N�mۦ���h{d�h۷o�B,����CH"����(Nj�Q� ��[�����C�P��� �)2����O�6�O�y.�7n���?����dB�s6m�dV�#gD��iDs/� |�5N� mp���?�X�	�H��H��hml�W�%�)Hf��xB��8+چI��G3P����G�82��h��?���_t$�|v��Q��'_�+d�4��×�7���*OM^uE�>N����ϟ_��6���iW�sZ�ɴ
������2�F��8X�bE�ş�]�v��T�
M"h��~�mi{\-O������[���?/���f���K�AM�;{Y$9�dR׮]]RM>��s	H��轗�э��ˇ�Xu�ƍt��ŧN�U�˄��J@4��[������)���.4Pwc$#++�5�\i*�W%�ߦ�ܹsG���I�n�@
};@῿��[�FO�P�(�T1@t���`4�zd��e��eV�.vKIe�J�����c'��kH��ɓ��菡n���;�y)���6c#�����Yg.�;��wlK�E&������ih⃶S�v�+  2��}���X
e,~�&���
�ՃS�q�i. L [�zɉD^��Cs`f�� u"`��ի�G���7�$2f��k���ccV�Z�ћ�{Bԙ3gʘ���4�z���[}���j��d<��b,@�7o^	 ��r��5ަ��_�Lc�Ȧ�:���Tho�ܨ�c�m�ܹ����'�,��>�Re1�ſ������ξ:\��L�Y�hQ1 ��(�Z��v>��j ��5;�ݻ����G�I@�È(  C֯_�˹��K�39 ����~.۱c�c���ݣ���%�I,^��dϞ=�� .�#&���� ��  ��/ƀ��nݺ�W�X�ޑ�ٳg%&����Z���dl�b!j_	ʯ�=veOb#��-Z���ꫯƶj��W|T�b<���T�^�Zb�@��ʟ�5�M�0a6�⢌���ѣG�5f������_$+�ѵ+s5r��o��@�KOOo�V�NHH���s��u���_<��̃�73aT�x�_!�A֐l0���`"*��<5}��X���GA�+���R��e�J	�߂�%����d��A ̳Os4����|���?~|�!�⓲�Ո�,���g�e&����55jT"+����9`� SZZZT����4_���B��K|�/�����l�_C��F ҋ`e՗ �)))�Æ����ɀdX]�?+�d�	8B�8�h�_#oC���8i& �<��7�z���}��c���$��Gc'k:�	��ը�w-c����h	��ԴiӐ�����#'�>�߯%�W����/� @8k@~��K��\ŚO��P��@W�&4D?�{��KKGS��޽{�F�t3۶m���X���.��%��ӌK���	�=j/�W�	6P�׼W�r
DXH@�������0���=���%̋0�ؤ��N�y��lOw��}�?b�ɶqX� �&���kf��Rܹ<�by��Q�����?��;���Y�������n�����LA[t�+�N��TX2�� &�{� �M"g�B���%M��b�Ii~��),���'K�Ÿsz��5mF�t �O�h��E�I�ND3�9K��\�CI�qI�� ��(�h�s�    IEND�B`�   g�8     8 �����8 (   O R   J u n c t i o n   ( o b j e c t )           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�[[[�ZZZ�ZZZ�^^^�___�^^^�YYY�ZZZ�\\\�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������nnn�eee�����������������������������bbb�uuu�����������������������������������������jjj�]]]�]]]�����������������������������aaa�����������������������������������������������������bbb���������������������������������lll�]]]�]]]���������������������ppp�����������������������������������������������������������������~~~�yyy�������������������������mmm�]]]�]]]�����������������bbb�����������������������������������������������������������������������������UUU���������������������nnn�]]]�]]]�������������UUU�������������������������������������������������������������������������������������ZZZ�����������������ooo�]]]�]]]���������ccc���������������������������������������������������������������������������������������������hhh�������������ppp�]]]�]]]�����yyy�����������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�����yyy�����������������������������������������������������������������������������������������������������hhh���������sss�]]]�\\\�kkk�������������������������������������������������������������������������������������������������������������xxx�����uuu�]]]�ZZZ�zzz�����������������������������������������SSS�111�111�111�111�333���������������������������������������������eee�����vvv�]]]�^^^�����������������������������������������777�111�PPP���������www�555�111�\\\���������������������������������������������www�]]]�[[[�������������������������������������LLL�111�uuu���������������������AAA�111�����������������������������������������ppp�www�]]]�^^^�������������������������������������111�???�����������������������������111�@@@�������������������������������������YYY�yyy�]]]�uuu���������������������������������uuu�111���������������������������������===�111�������������������������������������fff�uuu�]]]�~~~���������������������������������XXX�111���������������������������������[[[�111�������������������������������������nnn�ttt�]]]�������������������������������������;;;�111���������������������������������rrr�111�������������������������������������rrr�ttt�]]]�xxx���������������������������������???�111���������������������������������rrr�111�������������������������������������jjj�www�]]]�bbb���������������������������������[[[�111���������������������������������YYY�111�������������������������������������XXX�}}}�]]]�YYY���������������������������������xxx�111���������������������������������999�111�������������������������������������iii�~~~�]]]�___�������������������������������������111�888�����������������������������111�JJJ���������������������������������������������]]]�YYY�������������������������������������XXX�111�[[[���������������������666�111�������������������������������������rrr���������]]]�\\\�___�������������������������������������CCC�111�<<<�jjj��WWW�111�111�xxx�������������������������������������nnn���������]]]�]]]���������������������������������������������ppp�888�111�111�111�FFF�����������������������������������������}}}�������������]]]�]]]�����eee�����������������������������������������������������������������������������������������������������xxx�������������]]]�]]]���������ddd���������������������������������������������������������������������������������������������bbb�����������������]]]�]]]�������������```�������������������������������������������������������������������������������������UUU���������������������]]]�]]]�����������������UUU�����������������������������������������������������������������������������eee�������������������������]]]�]]]���������������������bbb���������������������������������������������������������������������ddd�����������������������������]]]�]]]�������������������������|||�qqq�����������������������������������������������������jjj�������������������������������������]]]�]]]���������������������������������sss�___�������������������������������������]]]���������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�rrr�jjj�ggg�eee�aaa�^^^�bbb�fff�iii�ppp�|||���������������������������������������������]]]�f% ;   % ��������G# �����$ /# ���������" ��������& �    O R   J u n c t i o n   ( o b j e c t ) 8   O R   J u n c t i o n   ( o b j e c t ) [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] 5 ����C p�  �����V@ �����V@          VUUUe/�@ ����ZR�@    �� J          �?�����F@�� J          �?�����F@ i             �����V@        �����V@ j5  ���� ���� � �          �! �����! �  ��������pL  �� K            S�����V@�� K            S�����V@         �� J          �?�����F@�� J          �?�����F@    �!  J          �?�����F@�C  J          �?�����F@ ib  �`  @   ~   ����?9@�����=P@�����'@������S@     q�      �        ��% % %                   r�                                            O s!     @@   @@   @@   @@ �       �B      �!                       {^!                          �^!       |�!                                       %�! �����!  ��!     ��!               ��!             ������!    O R   j u n c t i o n 9E" ����E" (   O R   J u n c t i o n   ( o b j e c t )         �8"     �E"        <S" ����S"  =�" �����"                       �?      �?                ?�" �����"  C�" ��������                              �?        t�"          ��U U U          �?u#   ��  ��� � �         u/#   ��    ��                                   m�$      n�# �t# k                ��# k          �?�����F@nF$ ��# j       �����V@��# j          �?�����F@��# j          �?�����F@�$ j                       �?         ݕk��|�?X���x�?n�$ �c$ b                  ��$ b          �����F@��$ j          �?�����F@��$ j       �����V@       �?         ӕk��|�?Y���x�?&% ��������2       �8 u  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�{pTE�o2Ʉ�x�@ !h�Ĉ��%�@�@�Ȣ��R�XP�]Y��t�c�(*B%�`�����G���Eނ<I&�d���ԝa&�sӷjj�ow�s~���ӧ�E�����J��y0nܸx��н���shhh\ccc\xxx;Σ��
		1𬺾��į�痸.�٥�����/_>�aÆ*=�I7 3fL,�MAx����Eh�&��KDDDm�����i�&�m۶111� ���]����(\�KJJjJKKk�^�Zw���Ѥ+7��IW�oyo���/�0��>���/6-22rBY]]�Э[7�m���������t��YAx�
͠ ��ɓʩS��9R~������� ����,m�(�{TP _*�1":66v�'��������Ԙ�}�����_���P:�V�ܹ3�rKjkk�VUU�^�z����r���CQ�ϡ��իWMZZZ��[���������ǕM�6��Ŷ���x-�	��+�0͂ u����ʝ Z?����?TK��'�!���+����h��`�d�������@���������ӧ��uL�޽�'�ʯ��P֭[W��W_Ր�n��\��g�2��K��h����f���t����?>�S�N>$�Y��ǖ-[?��S��_������W��K�B222G�;`����'F�E�֬�VP�94._��D�f��L��3���}P�'ӧ��رc�3bn������ʪU�j�����g��p��26�ݻ,��駟�2dH(�@�x�r����ŋW=z�<MD&�(
De��y�~�Z�Z����񩧞�ƃ�5UfAAAcvvv%��;h�4����_A@{?�nִi�"�*,����ʢE�*�L�ǐN��9~�������?mΜ917�t����r���B]NN�	��xz?�� �� I `۠A��_y����u�A�������2���)wx�޽{7�� ��  ��S��Ot���4���]��Th.�w�ؑB������s�ĉ_�3��KG��={v������]� ��
nr##���c<d���'�H��`D,��ʊ����]$_&o w@#�}/^�8���)x]#x�0D�C����o�3��D�����&M�nl,ƹԍ�C���Y��UM��AE�.\hA��h^CΜ9c@#���e���V�^��Q��`�cϞ=�U?�����sO@h˘C�=z�a#xũ���ޅ���y�u�W�kM�>��3�h�q�{��*�& �'#p۬Y�b����u�[��%�KHII	ߺuk� 
?�O���F�������;�Q^�Ғ����\ׯ_?��w?͂G��5�q�W+q���a-IZ�Ux^�ΝM��c�zz���KO`
���1�2����]�vah��.]���px�E�4������^���������h�	�{�|��w@�!��E+�r��>J>s��(���t�G�S�� �#���'F�l���a��΢�6.��� �&��s�ϟ/��]崏��|����z�ʕ���ٓ�Jq.i&�|��1�5��i1-��O�[��J����p�@����^���!|�Z�n��J�΂ ��&{���b��+�˴~���>
n��l�N��&`b|||ǁ:��L �譩S���N�etJ��(]·&O�,�$XW����;���.әw���R�s�w8��L�L�2%m�&�q8���, QRhD��VC��fl�5�Kw�N� (*:���R��Q��8��b�1��Qq͂ -0Wd�(�\�`)C��#��]�Xg���#2�Gpr@��9���<�9
삀�b����Ds��g��<�q?Q��WU� `M�i�����e(�k�"�0�zf5��W3� �G�l�R�����G�F���=6A@0�`�p{/����B��=HKOO���M0P�(�ʐ�����ڢ��k����Jtp.t5]�"m+��� L=��_mU�0�l��9�����+�	Y�4o �cB� 
^y۬9�)|�m����	n 	��R�u:y��u��<lM�p/��%lߵkW�t�Z��S�Y�b|��#��%�)h�=^w��=�A,�f$�2��ЂE���D�'�)k �(La���~�nA�X8�� ��8� �����|���&���5a �(L˧�C� �Ѐ��]M�x
x
�J�٣�sz~b� IM��-KO��;:<gN�����A  �G��b�:�eВ$��ad�����ׁ�#�Z� h9�+�&P�	,?3@G���ȗE22c1j�� �A}H	5wtx.���f�"�J�o��[�KaB�J��@� ��n}Q���Z
��E����ah�.�<�f�g	�C
��d�A��rFj�������V�&M�v�0�	�>8 v]������ڊKl�(�����sd}VM��W��Ds`%���\g`��z�]�CM��l`e��.���s�q����&��'�d�A�cx��U����8p�ܹz�j�,@@[q�������\g�t�pQ�eڊ�cǎU��s�p���T��vNM�N����K�9��s6����&��v��矑����i�u�s@l���������]�8�$#�q��_-c7��֔Y���Í���ѾJ�e�kp@hw��z�kQW6^�^ F��U�"�A��Z���4m� ��zQ Z�j�Νh����r֬Ys�����k+���ؾ}����U�@ 1漢������^�q���\9uꔈ+����M�4�lÆ�'�G��q�m�&&����l����	F��Y*ƚT���A�>�+�ګ�M����[��&r�e&�k��(Ǐc`0�^�� rvAAA(Ƅ�w�� � �j��5\�6�+H� �Iڑ�l���*��p}����D�-����]���`(oJ,���hrOxH�x�ռY�\�r=@8�k׮���4��W��^uT�fA ^���e$�k����S._�\��n����w��w�^mQ)k�,>���2�=/���\� �&�����ҥK�6h���y�8�B���}�L��@d����9Q�
��S�	 Ĕ��>��-��p�DU��ȌL�|���M�粉w�A�%l(++ۇX�l���B�q%ob�Q�)8�]?�E��y��4W�v"S�4}�Z�])C�����M4K�`]��]��U�N�^~���e0��$�d1�w�V0˙f6��W��\�����"�?���ܱw��.��\�<�*��(����	�m<���h w��H�3����f�#3s�hf�C��A#�ru
��I������[��;*C>�!~����C��a�X8��:\n�J9p��^���}�ȑ���w�\נ�1~�A?���	�<�o�q{&�� ��z����'��Q; �Q^~�.��M̟?s�bv�6O��Hph�z�T��I�S���#YA[.��4�|W�̛7� ��bŊl'_���#�\��TƖ9�1�<�o߾Ƹ�8����s@��.\hb����-[&\��@������i��Bw�]w�6+���*17�U�x��Y��-�ri�����-[��INNo׮�o�Ђs�0a�B/`n��X�E�)�Pѡ�҈��<����F�&O�\�����7�g��_l��G�~�m�ѣG�+[>s�D}+��e;v��CO�/��&@]�ךu�4�a,�ڼy�#��gd�M�cy�$D/��^�`L��������	� �@X�'��N��׵����db�~�rV[���o}6���~=�A7�G����;?�쳑���B�g�E��E�D ς���E�.�g����h�+����rV2�CW6m6��X�Ҕ��� A;uDp� �18�r����@�Z�,|�0�3-�/�III>�B�`�����eeeUǹ�Ć*�R`�'�� h��<��ӧO��ӧGK��lܸ�qɒ%�/D���@��h$~��@0���9�O�2%b���B5WO]>�HP�gp e���^������`���A�3f��z֥���1�Sj���Z� Y��=)
���	�l������Gdff�$$$X�Mר{�����J�-]�Y�b��@�\��&Bt�A1w�������(��A������/_.��v��Y;!p[ejM�1���0gS��ƈlzT�"�/_�ڵkk�����G �`��@�D�Q�"������1��HH���Y�F
ü
�
���>l����蟃Z��fA�f�  �B�>��6--�uJJ����p�k�lڴ���X4RX����,??���-��'���`*��N�:դ��F���/�G��?��;Ĉ5�Y$��a�0��s��~9���7������AÆk߾�O���n���F�-"�N*b��~��s�+b�w~|��D��Ju�:�25o_~����r�y!hA`�?�%�7�� ��!v'��ʿB�c��}��6m�D�I��rŞO�~��.�o�JJJ�q��b����	Gȑ���"�mBߊc�u��Z7 �'��c��!��|ѝ�Jv ]��܋�8�Y 0�w7�{��_D�'�?��/��l�^��}����r��r�e*+=��    IEND�B`�   g�d     �d �����d *   X O R   J u n c t i o n   ( o b j e c t )           �?�   !   !                                                                                                                               ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�\\\�ZZZ�[[[�___�ZZZ�UUU�ZZZ�UUU�[[[�```�ZZZ�[[[�\\\�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]���������������������������������hhh�www�������������������������������������mmm�ooo�������������������������������������jjj�]]]�]]]�������������������������jjj�������������������������������������������������������������uuu�����������������������������lll�]]]�]]]���������������������hhh���������������������������������������������������������������������aaa�������������������������mmm�]]]�]]]�����������������ZZZ�����������������������������������������������������������������������������UUU���������������������nnn�]]]�]]]�������������UUU�������������������������������������������������������������������������������������UUU�����������������ooo�]]]�]]]���������lll���������������������������������������������������������������������������������������������bbb�������������ppp�]]]�]]]�����bbb�����������������������������������������������������������������������������������������������������iii���������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�\\\�```�������������������������������������������������������������������������������������������������������������aaa�����uuu�]]]�ZZZ�������������������������������������555�111�������������������������AAA�111�������������������������������������{{{�����vvv�]]]�___�����������������������������������������111�GGG���������������������111�fff���������������������������������������������www�]]]�XXX�����������������������������������������KKK�111�����������������111�777���������������������������������������������ddd�www�]]]�eee���������������������������������������������111�444���������VVV�111�������������������������������������������������YYY�www�]]]�zzz���������������������������������������������ttt�111�ccc�����111�VVV�������������������������������������������������lll�ttt�]]]�����������������������������������������������������;;;�111�111�222�����������������������������������������������������sss�sss�]]]�}}}�����������������������������������������������������111�111���������������������������������������������������������mmm�uuu�]]]�qqq�����������������������������������������������������111�111�```�����������������������������������������������������ccc�xxx�]]]�\\\�������������������������������������������������333�777�999�111�����������������������������������������������������[[[�}}}�]]]�]]]���������������������������������������������XXX�111���������111�???�������������������������������������������������sss�~~~�]]]�]]]���������������������������������������������111�RRR���������XXX�111�|||�����������������������������������������������������]]]�[[[�nnn�������������������������������������999�111�����������������111�111�����������������������������������������aaa���������]]]�]]]�ppp���������������������������������iii�111�������������������������111�QQQ�������������������������������������������������]]]�]]]�����hhh�����������������������������111�AAA�������������������������AAA�111���������������������������������aaa�������������]]]�]]]��������������������������������������������������������������������������������������������������������������������������]]]�]]]���������ggg�����������������������������������������������������������������������������������������zzz�yyy�����������������]]]�]]]�������������WWW�������������������������������������������������������������������������������������UUU���������������������]]]�]]]�����������������eee�����������������������������������������������������������������������������vvv�������������������������]]]�]]]���������������������~~~�ppp�������������������������������������������������������������jjj���������������������������������]]]�]]]�����������������������������kkk����������������������������������������������uuu�ttt�������������������������������������]]]�]]]�������������������������������������zzz�[[[�sss���������������������ppp�___�������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�vvv�ooo�kkk�iii�hhh�kkk�ooo�vvv�~~~�������������������������������������������������]]]�faQ ;   aQ ���������O ����LQ �O ��������3O ��������' �    X O R   J u n c t i o n   ( o b j e c t ) 9   X O R   J u n c t i o n   ( o b j e c t ) [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] �K �����K pTK  �����V@ �����V@          VUUUe/�@ UUUUE��@    �)K J          �?�����F@�KK J          �?�����F@ i\K            �����V@        �����V@ j�K  ���� ���� � �          �{M �����M �L ��������p�L ��K K            S�����V@�
L K            S�����V@         �5L J          �?�����F@�WL J          �?�����F@    �}L J          �?�����F@��L J          �?�����F@ i�L ��L @   ~   �8��x�<@��8�C�N@�����'@������S@     qM     �        ��% % %                   rAM                                           X stM     @@   @@   @@   @@ �       �B      �{M                       {�M                          ��M       |�M                                       %�M ����LN  �N     �N               �+N             �����LN    X O R   j u n c t i o n 9�N �����N *   X O R   J u n c t i o n   ( o b j e c t )         ��N     ��N        <�N �����N  =�N �����N                       �?      �?                ?�N �����N  C3O ��������                              �?        tWO          ��U U U          �?uuO   ��  ��� � �         u�O   ��    ��                                   mLQ      n�O ��O k                ��O k          �?�����F@n�P �P j       �����V@�<P j          �?�����F@�^P j          �?�����F@�|P j                       �?         ݕk��|�?X���x�?nLQ ��P b                  ��P b          �����F@�Q j          �?�����F@�"Q j       �����V@       �?         ӕk��|�?Y���x�?&aQ ��������2       ��d i  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�	pU��o�"$�F�d	�����0$����:�*�T�࠭�ԥ:X,t�"j�2���E�� 6�&YdȒ�����1��ޗ�^�{y{Ν�s�s�9����~�;�wMS������V�x���۴i��7n$����R�谰�����r��x.)..��z��+�W�ބF��х
�߅�m[YYټ��<�����+�A-22�JN�� �ͳ��(��(�"�B@r����`EE�>��H}����9�a�G��J�fP�T^O*-�y��emڴ���;���[o�Ukܸ�+?��l� �v��y�~�������ĉ�˗/Ǒ�1�Z_RR�	��_�l���S�A�M�4����MEd6l�P�֭[��w������Un������k�}��y���׹����AB,ER,G�J���3f?ѝ���Vѿ�Į]�j͚5�[�O�fB;t萖��_�e˖*$��������Χ俘����&T��h�'%''G?��C{��v�-���cr�f������͛��m����d2���t���3�$Ǝ�N������3?������~g�+ 4�P�4@�(����*�ŢM�6�p%_�(P�ih�3h[�������>x5�={�h+W��v��I��+V����^�ԅ�T~�[�=~ذa�Ç�rV�w��~�*�CNNN�ٳg/�	�a�߉� � <;;�9�x���G>��#�� ���� �a޼y&��|�����G�7�9�c���hѢ�ĉ�y�^e|�%.]�5k�T.^����s�ν�/}�� @�GDGG���?���8p`x�U�/�cԜ9sL��"F �2�˧ ŏ�>755����?�ШQ#_�7`���`���J�;�aɒ%���P�� c�0 �	:@��H�*�,gP�UXX�͜9���ŋ[�
�
E� �56~��4��6mZ�]w��rm8��������]*++{  �va�
���-G����/6�>��+Ē�ƍ�}����cc�hy�k�7�4��{�m�m�ܹs��^z)!���❤��4�X̮]�Ƶk��6�����+ �>}>�ԧ�~:V���U�xD{���cǎA ����;�K��Wo�����~��#FD9�^�:��FN�4Iê��8�+q<*	�6E��!(D�B��k�bE0`��nݺ!;v,g�v��]� ���}��i��Ox,]׋�_0rJã�u��>4Wh�멒z��P�1���i T�ڱJG�лw�(���[�.@Y�u�&�p������#mܸq�Vt�Gs@�ŗ_~9���Hߞ�H�Β C�,�3ñ$�^�'���4�܎$�ڹs��V�Z}r�ȑk�e?F�@�)x���������WBd5?]����3�>�e�t7#��DQ;IӧO�����=�Eu��A�rs뒻[ ���bؿqǵlٲ.��o�ȁ�{N�_�%�r7)�@о}�L�h>x��:5'����?���S��#"�o���w.�@4R�L�<yr�s��~�ٶm[���9��� �EO=�T
�;��o���5��I��Ѯf��B_u�����q������F0AG�2e���>��1��� � ]�?�T"�1O���@c�VlRRҫ��45��̌���?W
W�J��rO��{���w
(���ÔY�Y��/�XQ���9�Y*�������&v6]Ϗ@'7�@����� Tuc!��4�&�G ʡ��at�Lgȩ����X�>�<4hP3������j� �G����<����q2�¥閙�X��F�C�����4���� �|���h�Qo|�:O �G	����xw����sD�]��H���o���� 
}M�dG%�F�>K����QF*�?`�Fs��d�a�� �6�yp� J�}��d: s>j�d� @�ݥK�
+��N�"���B/o�d� ���(�*G�=��{&k�{���w�Ez`r�an|/&�ڊ��)��~Cm�_(���J^"�:@���N��*QН�LX���V�cT������_��g�A���A\�H�w�����Vc֒b%dm�tF�JG�r����K�ߺ�5���%�TG�q 	�^�a]2쌩X5�\
�g6�XD��uq @�`���O`ͥyF'�X'1	���� �gЕ�N"�n]�����C��g :A�����&L=�����<M���#S��XϞл����E�Ʃ7¬X�z�W����`3h���� �B��C�������U����M�4��څ>Qu��!g(���b�   .��2�p��:6�1P���Qu=���M��I]�)4�@��mHc
0�'�E$J�6d�p)��5Pt,��f���k��c�^Y����_�+��]��.l��\_�j�,�AI=wB���ꋦ��k׮U?�#���� u,���/Qu���֭�AQ݇ؼ[c�y��4Ջ0��"���렏��C���
G�}i�%�g�}V,
Õ+W���>�8p�̙: '�Ū��ıpN��QG�r�=��i�O�Kh �?(��z��*u~\_2L&��'O�T�D=�B�^E4�2�쨾X�5�;z��O�����}Á�Q�*���w?������7�\|�u��u^�
_�b���
���g�x�98p��A��x�uQ �@��/+Y�S�!�@P�y�uQj� �p�*�YGT����^�~=i��$5@���˯����e��H=�����0[S_+W��#��.X�U�Á���"��r[E�"U�CX�g��V�ű |G�@ۻwov�/l�o���ꫯ���@�>|��2��ħ�~z���^D} �n�����|���V*� u�`��b#���6%��ݻ+��jǎ˒�D���倌$ڵkW�����	�L��.�eY�FÁ��<F��^S E���˗�!B~>|�p�@����_�v��]��&�F(�R�bI|�O����x��"8�����S6G,�0l>Ř��޴i�GT:��u�L|�>��0D�Q�*,08 N@D�P���(r��`����������%KJ0�c���ڨ������wSҠ6nH�ܶm[J�p��ZA ����3�J�8�R��Y�hQ1T�Ï��v
H�K(o̟?_��_�)`x�&^`���$�$"
�_lbڿ�<�#@9����a�=R���i�h9��fΜ9&ښ eA�&��/�4c8���_�p�iH� a5�վZ�x�y�
�}Wzo999e��~Mv.p	R2��v��2<�>(���Y̝;��m6?�!g���sdR�4xrƌ&��t�Տ৬,((8u���?�C�[S�q*f��t[���3ʝ��7�� L�Y�f�����YtѝT]��L�v��y�H5.Z⨫w9��F{���EQ	m�Z�J�n��Le����?���~p%O��q��g�.�a"ΩK�n�@2ňT���o�Ԭ��T���J=�������/��	�I0Q�HzzzV�>����s�;��ׯ7c���}�L�Q�5u�$|�����m۶F45�ԩS<#[���בLа
^C�I|������# ����۪�B2�`��hOT�1�~��<�#���?y�5C�8ۧN�*c�O����-]�T�ui�ԈP��BR���hi�C2�ѯ_?%�P9�O�	�`b�~ �e��%{W����	@X���ڙ�M���twK���ȁ�7��{�kH� ����NE�
�Y$�-[&S���vE�q��9�E��_�z͇�-�,-M�:�]��j�*J���'��/f�H��� '��ҽX^��D�q7:�vL�#�1DȎ�Yt��z�Uaa�6m�4өS�r��̡��{��>��Q�F������
m�L��Ш�ao�1h�fT�Y����&�,��^����x,B",`��5k�����Ql�h	��WYy��w�11��4
�@�2k}��I}��
�����:4~�g����~˖-U,(�!4?� ��K�R�C��INN~��������Lك�� @�	R�E� {s{��@�0�o �9r���l�8��6�M�0!�[�n����^�zU�j���@��Ο??�����f��A`)��ѣ�bK�Ӵi�&�?�xCQ�����r���
fF�����իWĪ�KM�;6�0���ј1c���[6n��Ufm��+ݼys]�%���#	�RA��a�!���'�A_�0`@d���$�~��Ϙ��_��G����w.�*�BK���B�FO�;�ĳ����۷�`�J���+�uW�	��cǎi۷o/�BZN��͢�1�_��� �p.+++G�HNOҕ� � Cb��ݵf͚Y���
0�"���-����M�ˡ��E�����!�����4��Is1
�?�T�`��2� --M�%K��?��=f\M�v��
�"b�`~��g�h��z$#'� ��=�t����b a��'6oܸq1ɪ���X�1<ktEo������,W #���b�M^N�2ssV����+\�������"�v�Z�*��	X�"###��f[޷cjVK$E;*/��<'Q�	\��{#9�����B���2���>��8�� �A�v�&wXӧ��������
    IEND�B`�	   g�     � ������     C o n n e c t i n g   a r r o w           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�����������������������������������������������������|||�����������������������������������������������������������������zzz�]]]�WWW�����������������������������������������������������ggg�XXX�nnn���������������������������������������������������������hhh�\\\�WWW�����������������������������������������������������fff�XXX�mmm���������������������������������������������������������hhh�\\\�]]]�����������������������������������������������������yyy�����������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�} ;   �} ���������| �����} y| ��������| ��������( �    C o n n e c t i n g   a r r o w 4   C o n n e c t i n g   a r r o w [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] sx �����x p6x �2w K    
   STUUU��u@         �qw K    -DT�!	@   
 <        ��w J   
        �?    (��@��w J           �?����*n�@    ��w J          �?TUUU��e@�	x J          �?         UUUUU�@ ����*n�@ UUUU�3�@ ����*n�@i>x            TUUU��u@                jsx  ���� ���� � �          �gz �����z �y ��������p�y ��x C   *   W      @��x C   *    X     �B@�y J    �'DT�!�? �'DT�!�? g        �-y J          �?TUUU��e@�Ey B         �B�    �ky J          �?      @��y J          �?     �2@ i�y ��y @   ~         @      @      @     `A@     q�y      �        ��% % %                   r/z                                             s`z     @@   @@   @@   @@ �       �B      �gz                       {�z                          ��z       |�z                                       %�z ����@{  ��z     �{               �{             �����@{    c o n n e c t i n g   a r r o w 9�{ �����{     C o n n e c t i n g   a r r o w         ��{     ��{        <�{ �����{  =�{ �����{                       �?      �?                ?�{ �����{  C| ��������                              �?        tA|          ��U U U          �?u_|   ��  ��� � �         uy|   ��    ��          ��| F                               m�}       n�| ��| j       TUUU��u@��| j          �?        nB} �} j                    �:} j          �?        n�} �b} j                    ��} j          �?        n�} ��} j          �?TUUU��e@��} j          �?        &�} ��������2       �� �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  aIDATx�رN�@`ۚ0��8���n��� �������d|	���	��q&�U�X$�z�@b@4���R��������Ύ @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� ���=��h4N�4=���N����/���`���lv�(�/
�jus��1�m��o̯��=V*��$In���]����u�r�\�`z�����&� sO�9��K����a&�y����Mx{��ڜ�_a�����}E_f��}����>A�һY�t4E��pa)\*���8�
�G������W�U,�n�;��f�2�Z�vp=�L[��Ӳ��-w!��x�*��iKnB  �������dvU0+;�8�6�*��n?��	 @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� ~.�7^�g�no�    IEND�B`�
   g�     � �����    C o n n e c t i n g   l i n e           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������|||�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f
� <   Ř ����Ř �� ��������Q� ��������� �    C o n n e c t i n g   l i n e 3   C o n n e c t i n g   l i n e [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] ~� ������ pA� �7� K    
   S��8�u@         �v� K    n���!	@   
 <        ��� B   
     %   ��8��Ɖ@�̓ B        %        0�@    �� J          �?��8�e@�� J          �?              P�@      0�@ �q�=�@      0�@iI�          ���8�u@      �      @j~�  ���� ���� � �          �o� ����� ֕ ��������p�� ��� E   *   ���8�u@�� M   *    X     �I@�� H    �'DT�!�? �'DT�!�? g        �/� H     Z��8�e@�M� H     [      �9�    �s� H          �?��8�e@��� I          �?     �9@ i�� ��� @   ~   ��8�e@��8�e@      $@     �D@     q�      �        ��% % %                   r7�                                             sh�      A    A    A    A �       �B      �o�      ��� ��� H          �?��8�e@                         {ޖ                           �ޖ       |�                                       %� ����v�  �&�     �:�               �O�             �����v�    c o n n e c t i n g   l i n e 9× ����×    C o n n e c t i n g   l i n e         ���     �×        <ї ����ї  =� �����                       �?      �?                ?� �����  CQ� ��������                              �?        tu�          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                 :
� ��������                                                        �� �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  :IDATx��1    �Om�@a��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`�<0� ���b    IEND�B`�   g��     �� ������ :   T e m p o r a l   I n d e t e r m i n a c y   M a r k e r           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�\\\�[[[�ZZZ�YYY�YYY�YYY�ZZZ�\\\�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]���������������������������������������������]]]�uuu���������������������ggg�kkk�����������������������������������������jjj�]]]�]]]���������������������������������ooo�}}}���������������������������������������������ddd���������������������������������lll�]]]�]]]�����������������������������ooo�������������������������������������������������������������aaa�������������������������mmm�]]]�]]]���������������������lll�������������������������������������������������������������������������fff���������������������nnn�]]]�]]]�����������������UUU���������������������������������������������������������������������������������eee�����������������ooo�]]]�]]]�������������sss�����������������������������������������������������������������������������������������vvv�������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������bbb���������rrr�]]]�]]]���������bbb�����������������������������������������������������������������������������������������������������www�����sss�]]]�]]]�����������������������������������������������������������������������������������������������������������������kkk�����uuu�]]]�]]]�����___�������������������������������������������������������������������������������������������������������������|||�vvv�]]]�]]]���������������������������������������������������������������������������������������������������������������������\\\�uuu�]]]�]]]���������������������������������������������������������������������������������������������������������������������{{{�mmm�]]]�]]]�lll���������������������������������������������������������������������������������������������������������������������hhh�]]]�\\\�YYY���������������������������������������������������������������������������������������������������������������������hhh�]]]�\\\�YYY���������������������������������������������������������������������������������������������������������������������iii�]]]�\\\�VVV���������������������������������������������������������������������������������������������������������������������iii�]]]�]]]�[[[���������������������������������������������������������������������������������������������������������������������iii�]]]�]]]�nnn���������������������������������������������������������������������������������������������������������������������lll�]]]�]]]���������������������������������������������������������������������������������������������������������������������ooo�uuu�]]]�]]]���������������������������������������������������������������������������������������������������������������������^^^��]]]�]]]�����___���������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������ccc���������]]]�]]]���������```�����������������������������������������������������������������������������������������������������������������]]]�]]]�������������ttt���������������������������������������������������������������������������������������������fff�������������]]]�]]]���������������������������������������������������������������������������������������������������������UUU�����������������]]]�]]]�����������������nnn�UUU�����������������������������������������������������������������������������XXX���������������������]]]�]]]����������������������www���������������������������������������������������������������������ccc�������������������������]]]�]]]�����������������������������aaa�������������������������������������������������������������ppp�����������������������������]]]�]]]�������������������������������������bbb������������������������������������������fff�������������������������������������]]]�]]]���������������������������������������������vvv�[[[�fff�rrr�zzz�qqq�[[[�ccc�������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�www�ttt�sss�rrr�uuu�{{{��������������������������������������������������]]]�f%� ;   %� ��������k� ����� S� ���������� ��������, �    T e m p o r a l   I n d e t e r m i n a c y   M a r k e r A   T e m p o r a l   I n d e t e r m i n a c y   M a r k e r [ I D E F 3   o b j e c t   s c h e m a t i c   s y m b o l s . c d l ] %� ����3� p�  ������H@ ������H@          ������@ �����o�@    ��� J          �?������8@�߭ J          �?������8@ i�            ������H@        ������H@ j%�  ���� ���� � �          �� ����}� t� ��������p<� �t� K            S������H@��� K            S������H@         �ɮ J          �?������8@�� J          �?������8@    �� J          �?������8@�3� J          �?������8@ iR� �P� @   ~   ������8@������8@������@���OUG@     q��      �      
  ��% % %                   rկ                                             s�                       �       �B      ��                       {L�                          �L�       |}�                                       %�� ���� �  ���     ���               ���             ����� �    t e m p o r a l   i n d e t e r m i n a c y   m a r k e r 9i� ����i� :   T e m p o r a l   I n d e t e r m i n a c y   M a r k e r         �\�     �i�        <w� ����w�  =�� ������                       �?      �?                ?± ����±  C�� ��������                              �?        t�          ��U U U          �?u9�   ��  ��� � �         uS�   ��    ��                                   m�      n² ��� k                ��� k          �?������8@nj� �޲ j       ������H@� � j          �?������8@�"� j          �?������8@�@� j                       �?         ݕk��|�?X���x�?n� ��� b                  ��� b          ������8@�ȳ j          �?������8@�� j       ������H@       �?         ӕk��|�?Y���x�?&%� ��������2       ��� l  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�]	pE��4�$�pDD 	�-.*^  ^`���W����Tai�Ȯl��,Rŵō�!� ��"f�<"�r$\!�~_�:5�|�޼{��]���������w����Bh�9�9�9`\h,���+k_z饙�ifԪU+�_���!<s���*��f͚�'O��X�z�	ħ�KY�|�͗Ԯ]��F�hG�0�!�<<7�s��>�������HJ�VTTl_�~�Y<{څ��6��[ni�7�:�/��'��Ћ�͋.�Ȁ�u���'=�+Ξ=+~��QYY)~��'�O�>��r|�7��b�}�ȑ#�
O�`ذa�!�� �� �VIկ_����3rss}NN�hڴ�����cM�8t��{��{��eee����y�m�@,A+-ZD�z�9�1�9��pv��0�ީS'^�k�N
>\a����'N�_}��رc�غu�طo�5�)й3/^�>���?���୿B�z0�&����&z��!=O��LW^^.JJJĦM��Ν;MТ�[��i?���U�VM&���VD��q5���B��/$A��ݻw7 :v��jg�p4�?�P�]�Vv#�:+�f����t���S��ɮ������9ޞ�7n�X\��b�����/�k���!tQZZ*V�\)���I��0후q�o�n��@�7�'��|72���[o�U\u�UIW��'�%4 ���$�9��t���)�U�NA���I^׀ ��c��������&����{^��� ,X �����E<�d�$�\h��h�T�>�n2�"�ի�p�$��m۶��3g���^V��`�3g]�|��DґT@ؙ�4�f6���@�3Fv�dB2�k֬���3���(�r��>L+�N]IT�������64��^�����8�|�7� �< �!��D�������m�q�W�GyDdff^��n7/�X%�Νk�|M�l�	{زe�ʪ��!� 4hPCx�C 9���?ޖ�8�-�Er�0e�e�>��F`*�6^�J�[�
�������=���;v��9?�`M����D���'�N��?r�������y�WCC���:�-����}vv�x��g��.�6�ǸI�QfI�w����O���2]��۷��1uq4@' `�n޶m[1a���;!�$gL\#���Ϲ1 @h  pA*f.� �(� ��y������ԺukѲeKc���B �	��&V���w9 �h��ڵ�x�'D�:�ť]$hѢ����7>��L"�:t� |IY�y�t����9EEE �㴋������o�/4�i �8�R}���b� ��7�D�q��	 +��{n֬���]4�5�5�¬��hJ��&�bO-���AP�/S���#͋��V���l�/���u ��H˫i�@�������k0�59lРA�d:.<x��_���b��b�ni�1��TN�Ο��������9�@aa!��q�R#�'�Y΁q)콌1�y �j�^�A���]�9 ��Ν;���b�ԩS��4֍Ć5  ���uϞ=ŨQ���z]C5xnF8cݺu�!����#�ʪ8x�Ř�)��������A�:I�9@K,�d���fa|pQ8uD�P�x��65jN�:m9 Y�6mڰĖ0��-����$�_��.����]�8 �x���|P� 4C/��DTr'@З�A=p�����q;����ɮ�xG�u�ȟt�l�zhw�u����9���X�����Og��uBID ��	ޜ�[����{8�E���[4�/��a��n�!����=Z���l�{����`
�H(R�L�cQh�`�"T���$q���oW5?j�|�Id�9RU�Cr�/)G���"�#1,@����%b�G0[��Oq��q�׎*� �cAlؕ��]��+4oޜ�Ĺ��v�9
�>����t�bW��w�������i�A�],ra@��c�;����Ïsqq�L˗���d!��+����y��c����A@�#���0P����[��8�s @f�B;�q�SEm���%t�oAH����W��`&�h�=p�Q���,��� $P� d�렡7����;��MgI,@�Y���� P�8��λ���C�^���%֖�`�l�λ�  �a W[[��8Yn�a��� ��֖��2172"�5�~� �%8/Gz�ȃ@27A�&|Gh��#�A5��Ĳp6@�:�k���P�׆���o���  b
�Pn`�.58`y��l�*[�6�ds���t+��2�W��d��V� ��ٗ"��}.O=؂ }F+&�Z@�*5B%O�Z�ق �"��xg�v�Á&M���@�K��-�)}��]�p�raH��m %�MׇLS l	![��fc߾Q{M@��L�KpY'Ȁ���򣒶� H��f'����`��Z�d�PZmA �e��]���D��IAh���4@kDS����m��{���08���}��` �	,TFz�����An�8+.L�1௖)�c�2����M�>^��� �kX`���-�/؂ 	+�R��\H��	� �˖ق F��Lp��Qڥ,�<��d$�����\�V�)�%Ot�e�9� �}|2*�S�J���|�$[�B�c�78;8r�W�i�
ؿ�l4�n�[0�2T:�Y;os�"����4�Lhɨ��Ѓ���~�+��oWM�-L���_��:�0���[���`'��=���&3!n�T�u�a(9���rUM	
��k���������*�=�^�C�:������-�Ox��Ν_~�%�𯷶!�&�eX�w�Z��g�q�]�I�����{���fضm�����&�l�c|�ƿ!A�t��чl���2,������cYRY.�'5$�}�B�7nd���8�)�o���ŋ�O�#�X��}����h�Ł�>�H�rp�":��o����,*6l����.� �q����@�:3��4���Bt�͛7���JZ	?Ŭ`k �� ��e(��pk��t�9��;�(�����1��3�^e˗/�/G�v!��~��7��pyy�\;��`o�kNa�h�ݻ׮L�`,')��JOۑV�XQ��Da�r�hW��O2v�ޭ��'a�܎��@�B0@���fYY��s!,X��z�/��(>"�c��ف��qI��֭[Ei��vv�)��	,���())	U��?��j�Y�d�躟_�jU�3���[x�5�B���@)��j��Ղ�I�ݘͽ"��;"0gEE�4TTJ��$:au��P��ϗ�A��qN��1x���>Trn�ʕ&��i�\L�>�Z����K�,����*b�`KP�?��_��B(n���5k���_�G���SUT `E�D�G�����-���إݷo��3g�Z$��[o�uv0j����w�IU����s;�:*�'ĦN��/�p���X�(�%Q� `Y@�������^�&e2"A���_���aWxX݀"��z�6ܱcGI�Z�?*���w=k����A8�1��X ��~����̓d��_1��R���-/����蕅1�~,..V�A(��wC��i��˳�gg���!��D��ݹG1R�t� ��� ��2��'�fH�8*� `��N�k��} �N�U�x�[�n�E<�]��/�`��/� �\����9X%�;��`Gb'R�cǎ�.]�h ��G��5<q�D3�fA<4��?�֍�a��O�n�5�6M��kYw%㗌�� �" ��� N~��/i�?�R�����܇S#p����5�Zm�Lp{��N�<�'��� �(t��@L\BFl���;4�4��i�F�7N���Ť�^7�b��7	�i�B�c���JB#�F�n����Z��M�na����q�_y��7�>CC��	 �8$S�a���LH��
 a�`�KK��M����ˋ��͉�5g ��O?eO�  ���0�z �g a31���FҖPPP �7���Jʃ��&M2<Ȯ���k�ދg2&Ԁ�Ç����.�F���⡇;v���)!�KR�o�J� 0 �����1�A�o�����W_-F�u�]�ţb3f�0aO�<NAK��B�n'�b������n윉����ޘB�Z�v���r��8�,)��{0^y����`�1 p#  ���ƺ��C�m��4�?ϋ���iiL3U-��c����C�C��C��b>��.׀@�.b8�'÷b\۶m�m���B�����q�˿�� ��BB�g�]6����p=�x;��oʸ��\���E�^�<wM�mb�_~' �}�������ml_2�+A�2hР����a�~`�a<��5���g8��x��M!�n���砾��C�4�����-���I�xG#�1r�T��oժ��=z����*:i!��=��N��~K�B�?���������Y��bO��J7�!�b�~č��^� �����������1}�!G~���M�{U	��~��Y�A`��w[XM��E��Sע��~0��z'�/c�f�D~~��ep<���#h�����'N�/����Z�"�@T��j��K@� d!f ߇j���,�� h���:��Dw��5�'�+7ṉ��u�ԑ� 8 *��zZ�xi�O[>U��ۅ��Q���뿛�Q�}!�S����VVV�EPD{t>|K�HdGQV��Dy� L)����#��.%A`'��I�&��S�2 �<ׇ����5�m&����9�yu�~�8B�444444444R����6�8,~    IEND�B`�   gC�     ?� ����L� ,   U n i t   o f   B e h a v i o r   ( U O B )           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�YYY�������������������������������������������������������������������������������������������������������������������������iii�]]]�����������������������������������������������������������������������������������������������������������������������������UUU�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������[[[�\\\�����������������������������������������������������������������������������������������������������������������������������YYY�\\\�������������������������������������������������������������WWW�������������������������������������������������������������UUU�[[[�������������������������������������������������������������___�������������������������������������������������������������ZZZ�[[[�������������������������������������������������������������___�������������������������������������������������������������ZZZ�[[[�������������������������������������������������������������___�������������������������������������������������������������ZZZ�[[[�sss�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�XXX�uuu�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�UUU�[[[�XXX�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f^� 5   ^� ��������V� ����V� � �    U n i t   o f   B e h a v i o r   ( U O B ) ;   U n i t   o f   B e h a v i o r   ( U O B ) [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] �� ������ p]�        |@      @o@               ]�@ VUUUu�@    �2� J          �?      l@�T� J          �?     @_@ ie�    
qV~B��      |@���e|�|�     @o@ j��  ���� ���� � �          ��� ������ �� ��������p�� ��� K            S      |@�� C        
ףp=g@         �6� J          �?      l@�T� J                    �z� J          �?      l@��� J                 i�� ��� @   ~   ��8���_@�q\-t@
ף�{Q@
ףȒ�\@     q	� 
    �        ��% % %                   r:� 
                                       
   U O B   L a b e l s s�     �A   �A   �A   �A �       �B      ���      ��� ��� J                ��� J                �� ��� J                �� J            @o@�M� �'� J             |@�E� J                ��� �h� J             |@��� J            @o@                {��                           ���       |��                                       %� ����m�  ��     �%�               �:�             �����m�    u n i t   o f   b e h a v i o r ,   U O B 9�� ������ ,   U n i t   o f   B e h a v i o r   ( U O B )         ���     ���        <�� ������  =� �����                       �?      �?                ?!� ����!�  CV� ��������                              �?        V� ��������A� ����A�    f}� ;   }� ������ � ����h� �� ���������� ���������            � ������ p�� ��� O	            S      |@�#� O	            S     @o@         �O� N          �?      l@�r� N          �?     @_@    ��� J          �?      l@��� J          �?     @_@ i�� ��� @   ~                 |@             @o@ j�  ���� ���� � �          �                     {\�                           �\�       |��                                        %�� ������  ���     ���               ���             �������     9� �����             ���     ��        <� �����  =P� ����P�                       �?      �?                ?^� ����^�  C�� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                    mh�      nZ� �4� k                �R� k                n�� �z� j    � ��D=��RB���=��� j            @o@n�� ��� j             |@��� j            @o@n$� ��� j             |@�� j                nh� �A� b                  �`� b                  &}� ��������2       f_� ;   _� ����h� �� ����J� �� ��������u� ���������            � ����� p�� ��� G          �?      l@�'� K	         Z�����?S�Q��IP@         �O� N                �n� N            @o@    ��� J                ��� J       �Q��IP@ i�� ��� A   ~                 l@        �Q��IP@ j�  ���� ���� � �          ��� ����o� R� ��������p� �R� K            S      l@�|� K            S�Q��IP@         ��� J          �?      \@��� J          �?�Q��I@@    ��� J          �?      \@�� J          �?�Q��I@@ i0� �.� @   ~   �q'i6@�q�Ri@�G�:��&@�Q�n��J@     q�� 
    �      
  ��% % %                   r�� 
                                       
   N o d e   R e f   # s��      A    A    A    A �       �B      ���                       {>�                           �>�       |o�                                        %}� ������  ���     ���               ���             �������     9�� ������             ���     ���        <�� ������  =2� ����2�                       �?      �?                ?@� ����@�  Cu� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                    mJ�      n<� �� k                �4� k                n�� �\� j    � ��D=��RB���=�z� j       �Q��IP@n�� ��� j             l@��� j       �Q��IP@n� ��� j             l@��� j                nJ� �#� b                  �B� b                  &_� ��������2       fA� ;   A� ���������� ����,� �� ��������W� ���������            �� ������ p�� ��� G          �?      l@�	� K	         Z�����?S�Q��IP@         �1� N             |@�P� N            @o@    �r� J             l@��� J       �Q��IP@ i�� ��� A   ~                 l@        �Q��IP@ j��  ���� ���� � �          ��� ����Q� 4� ��������p�� �4� K            S      l@�^� K            S�Q��IP@         ��� J          �?      \@��� J          �?�Q��I@@    ��� J          �?      \@��� J          �?�Q��I@@ i� �� @   ~   �8��(9@�8����h@�G�:��&@�Q�n��J@     qd� 
    �      
  ��% % %                   r�� 
                                       
   I D E F   R e f   # s��      A    A    A    A �       �B      ���                       { �                           � �       |Q�                                        %_� ������  �h�     �|�               ���             �������     9�� ������             ���     ���        <�� ������  =� �����                       �?      �?                ?"� ����"�  CW� ��������                              �?        t{�          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                    m,�      n� ��� k                �� k                nd� �>� j    � ��D=��RB���=�\� j       �Q��IP@n�� ��� j             l@��� j       �Q��IP@n�� ��� j             l@��� j                n,� �� b                  �$� b                  &A� ��������2       R� ��������       �^�   �?� �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  BIDATx�YlMk�W�C)5��1DW$�1FnBx �� 1{h"�"1�A�Ĕ��PS��)fAH̪B���������)=����[Y���9�{�}��o���}{��-�F$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@$@q$L�0�/oz��2J���8����
���s��5*���X�|yq�ڵ3B�j�*���L��}6	4k֬����hSU��	\h��	�&�EM�B�h,M`4�.�hZFci��u�E��2KM��,�����X��hb]d�.����F�"�&p�e4�&0�XY4�-��4��ĺȢ	\h��	�&�EM�B�h,M`4�.�hZFci��u�E��2KM��,�����X��hb]d�.����F�"�&p�e4�&0�XY4�-��4��ĺȢ	\h��	�&�EM�B�h,M`4�.�hZFci��u�E��2KM��,�����X��hb]d�.����F�"�&p�e4�&0�XY4�-��4��ĺ�
}��%��ɓ.ǘ�MLL�Y@�4STTBl����)7n�z���{��I^^����۔��b�?�ZRR���T2s�̄�Z�[�d��k�N�'�Y�X˓'O�����5A`dvi����&��n M`7����%B��'NH�*U�G�r��-	�BҪU�X�D�_�pAn޼hх�y���$%%I˖-�u�֑���ȑ#r���޽��1⇐k׮I�-�Ν;Ҷm[�V��1A6�<�=�Ќ�y���a�`P�~}�ԩ��A���?�����<x�ߤ�:t��M�F���U����`�ڵ2k�,��B��=*A�)�x�Bn߾��0.^�(S�L��۷���,^�X����k׮eƭY�F�V�*�{�A6ʖ-[�������G��͕;vȥK�d���2d�y����	`��ׯ����e�3��_�~]��q+zۭ[7ٰa������g�d�Ν:�.�5�ϟ?��͛5��M���ڵk�<|�P۹s��S�g$�K�.ұcG=ovv�xװr��ٿ�4n�X&N�(��}u$�>}Z��߿/x���;&�޽�s��鈌���gϞ�w�^eмys=�g����&��ɑݻw��cǎU��

�����7�b����g�z<n�8���=z�4h�@�W��������X�B+ŠA��N�:zc���Z� x87Fs��$���֭[�Ɇ�֯_/M�4�Z)5��#�1�PQ�g k?�����U�y��I�t�@�C۳g��Z�J_��006mڤ�x��(�?��S�e�ȑZ6l��0:۴i�F����W�ʡC�d�ҥ���Çr��)9��»1���4w��-5b�cѢE����9�p^��+W����
C]�|Y���1�`��g��1��P����jXk���	j֬)u��կ�N���_	ʺE]��j3f�:T��TLX���shzz��Y�����a�ԩ:RKy�L�6M���#S���O�Jrr���������"��
�4c4aQ�n�cp��0���.fq�~���2�?@�o���Q��:��(�(�~�ýv�F$�q���s5�7F,��#�}����|�S�^=�����̙�U�b���=�D��\�n�^�\�R�Ѷm��� 0ۼy�t��o�>��W��@&@gG���1�8PW�x!	X0a�֧O9|��$$$HZZ���ɓ'˰a��(F���h,��˖-,� {���ҿ=���E��8L���я��>�����̸j��̔ٳgG�0c�5;��^�V����oܸ����8�R\��r�oޯ�:z���˗/u�W���w��1=`���? ��w������W��RN�5A,�ы?&%%E�*��˲���V�F�x�M��?��L����h�Jn �O�xszIed���']Ur���{�iޫ���J���b�R�RVD��UѾ}��*Q�)�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H���ߒ�E�_{y�    IEND�B`�   gS     O ����\ ,   S i m p l e   P r e c e d e n c e   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������|||�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�fv <   1 ����1  ��������� ��������F �    S i m p l e   P r e c e d e n c e   L i n k ;   S i m p l e   P r e c e d e n c e   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] � ���� p� �� K    
   S    Ao@         �� K    n���!	@   
 <        �! B   
     %      @Pt@�L B        %        P�@    �r J          �?    A_@�� J          �?               i@      P�@    � |@      P�@i�          �    ao@      �      @j�  ���� ���� � �          �� ����_ V ��������p �@ E   *   �    Ao@�a M   *    X     �I@�� H    �'DT�!�? �'DT�!�? g        �� H     Z    A_@�� H     [      �9�    �� H          �?    A_@� I          �?     �9@ i4 �2 @   ~       A_@    A_@      $@     �D@     q�      �        ��% % %                   r�                                             s�      A    A    A    A �       �B      ��                       {.                           �.       |_                                       %m �����  �v     ��               ��             ������    s i m p l e   p r e c e d e n c e   l i n k 9/ ����/ ,   S i m p l e   P r e c e d e n c e   L i n k         �"     �/        <= ����=  =z ����z                       �?      �?                ?� �����  C� ��������                              �?        t�          ��U U U          �?u�   ��  ��� � �         u   ��    ��                                :v ��������                                                        �O �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  :IDATx��1    �Om�@a��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`�<0� ���b    IEND�B`�   g5;     1; ����>; D   G e n e r a l   C o n s t r a i n t   P r e c e d e n c e   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�����������������������������������������������������|||�UUU�UUU�UUU�����������������������������������������vvv�}}}�����zzz�]]]�UUU�bbb�ccc�ddd�ddd�ddd�ddd�ddd�ddd�ccc�ccc�ccc�ccc�ccc�YYY�UUU�UUU�UUU�aaa�ccc�ccc�ccc�ccc�ccc�ccc�ccc�ccc�ccc�___�UUU�UUU�fff�]]]�\\\�����������������������������������������������������www�UUU�UUU�UUU�����������������������������������������qqq�ddd�����{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�7 5   �7 ��������5. ����5. � N "   G e n e r a l   C o n s t r a i n t   P r e c e d e n c e   L i n k G   G e n e r a l   C o n s t r a i n t   P r e c e d e n c e   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] C* ����Q* p* �) K    
   S     @o@         �A) K    -DT�!	@   
 <        �i) J   
        �?WUUUUg�@��) J           �?    ؃@    ��) J          �?     @_@��) H          �?         WUUUU�@     ؃@ WUUUUO�@     ؃@i*                 @o@      .�        jC*  ���� ���� � �          �7, �����, �+ ��������pf+ ��* C   *   W      @��* C   *    X     �B@��* J    �'DT�!�? �'DT�!�? g        ��* J          �?     @_@�+ B         �B�    �;+ J          �?      @�]+ J          �?     �2@ i|+ �z+ @   ~         @      @      @     `A@     q�+      �        ��% % %                   r�+                                             s0,     @@   @@   @@   @@ �       �B      �7,                       {v,                          �v,       |�,                                       %�, ����4-  ��,     ��,               ��,             �����4- "   g e n e r a l   c o n s t r a i n t   p r e c e d e n c e   l i n k 9�- �����- D   G e n e r a l   C o n s t r a i n t   P r e c e d e n c e   L i n k         ��-     ��-        <�- �����-  =�- �����-                       �?      �?                ? . ���� .  C5. ��������                              �?        �7 ���������7 �����7    f�2 ;   �2 �����2 �1 ����p2 �1 ��������_1 ���������            �/ ����Y0 p�/ ��. K	            S     @o@�/ K	            S                 �./ J          �?     @_@�Q/ J          �?            �w/ J          �?     @_@��/ J          �?         i�/ ��/ @   ~                @o@                            �                     {(0                           �(0       |Y0                                       %g0 �����0  �p0     ��0               ��0             ������0     9�0 �����0             ��0     ��0        <�0 �����0  =1 ����1                       �?      �?                ?*1 ����*1  C_1 ��������                              �?        t�1          ��U U U          �?u�1   ��  ��U U U         u�1   ��    ��                                   mp2       n*2 � 2 j                �"2 j          �?        np2 �F2 j            @o@�h2 j          �?        &�2 ��������2       f�7 ;   �7 ��������K6 �����7 36 ���������5 ��������� L         4 �����4 p�3 �3 C         >@ |       >@�(3 C         >@ |       >@         �T3 J          �?     @_@�w3 N          �?            ��3 J          �?      .@��3 J          �?      .@ i�3                  >@              >@ j4  ���� ���� � �          �                     {R4                           �R4       |�4                                       %�4 �����4  ��4     ��4               ��4             ������4     9�4 �����4             ��4     ��4        <	5 ����	5  =F5 ����F5                       �?      �?                ?T5 ����T5  C�5 ��������                              �?        t�5 ��5 F                ��U U U          �?u	6   �� ��5 F   - ��U U U ��5 F           �6 F        u36   ��    ��  �+6 F                                        m�7      n�6 �x6 k                ��6 k                n�6 ��6 j                ��6 j             >@n"7 ��6 j             >@�7 j             >@nd7 �>7 j             >@�\7 j                n�7 ��7 b                  ��7 b                  &�7 ��������2       �7 ��������    L ��7   �1; N  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�ٿ�SA�f_�R�V;�F����И<��o`c'�bi�V�	DS���� *� h�O���Y�����aaNΜo~dsw��| @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @ +�d�R�����z�{��V�/���n�����`p�i�ϣ��M��~��+u��8���y�(S�r͕��p�"�>̄�L���?DX���"�#���T�Fj��|�0ܬ�l��f�W!�(w�f�0AG.�8��W�xĸ.�ɖמ��3~�߯ϒ����l��ѵ�f1�*�^�������~��)^�}͋tl��8{�E�l�ͅ��b���\����&��Um�.��s��{��璵���;�����6��8�͞L���f��XT=��/��A������_F�"�[�F�_F�"�k�嗑��Ht{M]~y�C����?�O��5k|��Z��$�.��W1���?��9�$@�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� �S)��9�����    IEND�B`�   g�_     �_ �����_ H   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�[[[�����������������������������������������������������jjj�bbb�������������������������������������������������YYY�jjj�����zzz�]]]�VVV�hhh�jjj�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�XXX�UUU�UUU�```�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�iii�WWW�UUU�[[[�nnn�]]]�]]]�����������������������������������������������������rrr�����������������������������������������������������ccc���������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�\ 5   �\ ��������+S ����+S � S $   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k I   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] 1O ����?O p�N ��M K    
   S     @o@         �/N K    n���!	@   
 <        �WN J   
        �?������@�N J           �?�������@    ��N J          �?     @_@��N J          �?         �����2�@ �������@ ������@ �������@i�N                 @o@      .�        j1O  ���� ���� � �          �%Q �����Q �P ��������pTP �sO C   *   W      @��O C   *    X     �B@��O J    �'DT�!�? �'DT�!�? g        ��O J          �?     @_@�P B         �B�    �)P J          �?      @�KP J          �?     �2@ ijP �hP @   ~         @      @      @     `A@     q�P      �        ��% % %                   r�P                                             sQ     @@   @@   @@   @@ �       �B      �%Q                       {dQ                          �dQ       |�Q                                       %�Q ����&R  ��Q     ��Q               ��Q             �����&R $   d i r e c t i o n   c o n s t r a i n t   p r e c e d e n c e   l i n k 9�R �����R H   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k         ��R     ��R        <�R �����R  =�R �����R                       �?      �?                ?�R �����R  C+S ��������                              �?        �\ ���������\ �����\    f�W ;   �W �����W �V ����yW �V ��������hV ���������            �T ����bU p�T ��S K	            S     @o@��S K	            S                 �$T J          �?     @_@�GT J          �?            �mT J          �?     @_@��T J          �?         i�T ��T @   ~                @o@���ư����ư> j�T  ���� ���� � �          �                     {1U                           �1U       |bU                                       %pU �����U  �yU     ��U               ��U             ������U     9�U �����U             ��U     ��U        <�U �����U  =%V ����%V                       �?      �?                ?3V ����3V  ChV ��������                              �?        t�V          ��U U U          �?u�V   ��  ��U U U         u�V   ��    ��                                   myW       n3W �	W j                �+W j          �?        nyW �OW j            @o@�qW j          �?        &�W ��������2       f�\ ;   �\ ��������T[ ����w\ <[ ���������Z ��������� L         Y �����Y p�X �X C         >@ |       >@�1X C         >@ |       >@         �]X J          �?     @_@��X N          �?            ��X J          �?      .@��X J          �?      .@ i�X    ���ư�      >@              >@ jY  ���� ���� � �          �                     {[Y                           �[Y       |�Y                                       %�Y �����Y  ��Y     ��Y               ��Y             ������Y     9Z ����Z             ��Y     �Z        <Z ����Z  =OZ ����OZ                       �?      �?                ?]Z ����]Z  C�Z ��������                              �?        t�Z ��Z F                ��U U U          �?u[   �� ��Z F   - ��U U U ��Z F           �[ F        u<[   ��    ��  �4[ F                                        mw\      n�[ ��[ k                ��[ k                n�[ ��[ j                ��[ j             >@n3\ �	\ j          �?      >@�+\ j          �?      .@nw\ �P\ b                  �o\ b                  &�\ ��������2       �\ ��������    L ��\   ��_ .  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�ؽn�P`'"׀�C7����!�W {/����&���*$����be ���
UD�=�:�d���|���rRU6 @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� 6L����������d2�짾i*t�b�ub���ç����l6{�kaHmw�/S�Ǯa("������]Cj{�5%���x	C#�~,1�0A����0�|%�L��I�a��Y��ʗ��xxUeW^��G��v�z~�V���9���s�mxj�˗�����)s^-�˷���y�,���@}���!���N��X7y���چ�<����.����l���]��x���%4������:,�<IC�l���;�~�X,~6s.�͋�{�����g�cAU�|!��&U�W������Ϳ���B�"w�_6����2����}���,�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� ���t��}�    IEND�B`�   g*�     &� ����3� Z   O p p o s i t e   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�[[[�������������������������������������������������������������YYY���������������������������������������������VVV���������{{{�]]]�VVV�hhh�jjj�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�jjj�\\\�UUU�UUU�^^^�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�aaa�UUU�UUU�nnn�yyy�]]]�]]]�������������������������������������������������������������zzz���������������������������������������������ppp���������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�� 5   �� ��������4x ����4x � T -   O p p o s i t e   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k R   O p p o s i t e   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] t ����$t p�s ��r K    
   S     @o@         �s K    n���!	@   
 <        �<s J   
        �?�q�qu�@�ds J           �?�����"�@    ��s J          �?     @_@��s J          �?         �q�q��@ �����"�@ �q�q]�@ �����"�@i�s                 @o@      .�        jt  ���� ���� � �          �
v ����zv qu ��������p9u �Xt C   *   W      @�yt C   *    X     �B@��t J    �'DT�!�? �'DT�!�? g        ��t J          �?     @_@��t B         �B�    �u J          �?      @�0u J          �?     �2@ iOu �Mu @   ~         @      @      @     `A@     q�u      �        ��% % %                   r�u                                             sv     @@   @@   @@   @@ �       �B      �
v                       {Iv                          �Iv       |zv                                       %�v ����w  ��v     ��v               ��v             �����w -   o p p o s i t e   d i r e c t i o n   c o n s t r a i n t   p r e c e d e n c e   l i n k 9�w �����w Z   O p p o s i t e   D i r e c t i o n   C o n s t r a i n t   P r e c e d e n c e   L i n k         ��w     ��w        <�w �����w  =�w �����w                       �?      �?                ?�w �����w  C4x ��������                              �?        �� ���������� ������    f�| ;   �| �����| �{ �����| �{ ��������q{ ���������            �y ����kz p�y ��x K	            S     @o@�y K	            S                 �-y J          �?     @_@�Py J          �?            �vy J          �?     @_@��y J          �?         i�y ��y @   ~                @o@                 j�y  ���� ���� � �          �                     {:z                           �:z       |kz                                       %yz �����z  ��z     ��z               ��z             ������z     9�z �����z             ��z     ��z        <�z �����z  =.{ ����.{                       �?      �?                ?<{ ����<{  Cq{ ��������                              �?        t�{          ��U U U          �?u�{   ��  ��U U U         u�{   ��    ��                                   m�|       n<| �| j                �4| j          �?        n�| �X| j            @o@�z| j          �?        &�| ��������2       f�� ;   �� ��������]� ����|� E� ��������� ��������� L         ~ �����~ p�} �} C         >@ |       >@�:} C         >@ |       >@         �f} J          �?     @_@��} N          �?            ��} J          �?      .@��} J          �?      .@ i�}                  >@              >@ j~  ���� ���� � �          �                     {d~                           �d~       |�~                                       %�~ �����~  ��~     ��~               ��~             ������~     9 ����             �      �        < ����  =X ����X                       �?      �?                ?f ����f  C� ��������                              �?        t� �� F                ��U U U          �?u�   �� �� F   - ��U U U �� F           �� F        uE�   ��    ��  �=� F                                        m|�      n�� ��� k             >@��� k                n� �̀ j             >@�� j             >@n8� �� j                �0� j          �?      .@n|� �U� b                >@�t� b                  &�� ��������2       �� ��������    L ���   �&� o  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx��1��p��Y�"�T
"��PD��cѩH���$���twrrpִ�~���p����p���$О"MM��ڴ���������� @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @������n2���v�w������;.�z�G�N�h�X|+R�~�EU_�?�d�Z5�;e��lD}����q�������+kb�Ï�����˥~�^��ABn��6�E�P�Ti��Z����/�Z��N�������W��.������VlW�^��q�{_b����~����/��i�$/����r�1N�&�v��h8������9��Ǘ�&z�}��I��6��.�ؙ�@i��?��Il7�9_ ��O��m�����v�����{�D?�b��f���l��7A�S���t:}}&yð�6�~�S�B��]�0�v�F]C��_�0l5���!���\�Ϛ�L���Oa�|��{��_�nJVX�k�z�j�('�J>?��m<i�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� ���6��͉�	`    IEND�B`�   g�     � ������ T   B o t h   D i r e c t i o n s   C o n s t r a i n t   P r e c e d e n c e   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]���������������������������������������������������������ggg�]]]���������������������������������������������������������zzz�]]]�YYY�����������������������������������������������������___�UUU�UUU�ZZZ�����������������������������������������XXX�YYY�����www�]]]�XXX�������������������������������������������������|||�WWW�UUU�UUU�UUU�ttt�������������������������������������XXX�UUU�lll�rrr�]]]�]]]���������������������������������������������������������ZZZ�VVV���������������������������������������������www���������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f� 5   � ��������\� ����\� � U *   B o t h   D i r e c t i o n s   C o n s t r a i n t   P r e c e d e n c e   L i n k O   B o t h   D i r e c t i o n s   C o n s t r a i n t   P r e c e d e n c e   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] J� ����X� p� �	� K    
   S    @o@         �H� K    n���!	@   
 <        �p� J   
        �?�������@��� J           �?:��8��@    ��� J          �?    @_@��� J          �?         �������@ :��8��@ �����y�@ :��8��@i�                @o@ H��65�        jJ�  ���� ���� � �          �>� ������ �� ��������pm� ��� C   *   W      @��� C   *    X     �B@�� J    �'DT�!�? �'DT�!�? g        �� J          �?    @_@�� B         �B�    �B� J          �?      @�d� J          �?     �2@ i�� ��� @   ~         @      @      @     `A@     q՚      �        ��% % %                   r�                                             s7�     @@   @@   @@   @@ �       �B      �>�                       {}�                          �}�       |��                                       %�� ����K�  �ś     �ٛ               ��             �����K� *   b o t h   d i r e c t i o n s   c o n s t r a i n t   p r e c e d e n c e   l i n k 9Μ ����Μ T   B o t h   D i r e c t i o n s   C o n s t r a i n t   P r e c e d e n c e   L i n k         ���     �Μ        <ܜ ����ܜ  =� �����                       �?      �?                ?'� ����'�  C\� ��������                              �?        � ��������ͦ ����ͦ    f�� ;   �� ����ȡ � ������ �� ���������� ���������            � ������ pɞ ��� K	            S    @o@�)� K	            S                 �U� J          �?    @_@�x� J          �?            ��� J          �?    @_@��� J          �?         i�� �ޞ @   ~               @o@                 j�  ���� ���� � �          �                     {b�                           �b�       |��                                       %�� ����ܟ  ���     ���               �ӟ             �����ܟ     9� �����             ���     ��        <� �����  =V� ����V�                       �?      �?                ?d� ����d�  C�� ��������                              �?        t��          ��U U U          �?u۠   ��  ��U U U         u��   ��    ��                                   m��       nd� �:� j                �\� j          �?        n�� ��� j           @o@��� j          �?        &�� ��������2       fͦ ;   ͦ ��������K� ������ 3� ���������� ��������� Y         � ������ pȢ   H��6E@  H��6E@         �T� J          �?    @_@�w� N          �?            ��� J          �? H��65@��� J          �? H��65@ iТ             H��6E@         H��6E@ j�  ���� ���� � �          �                     {R�                           �R�       |��                                       %�� ����̣  ���     ���               �ã             �����̣     9�� ������             ��     ���        <	� ����	�  =F� ����F�                       �?      �?                ?T� ����T�  C�� ��������                              �?        t�� ��� F                ��U U U          �?u	�   �� �פ F   - ��U U U �� F           �� F        u3�   ��    ��  �+� F                                        m��      n�� �|� k          �? H��65@��� k                n� ��� j                �� j          �? H��65@n.� �� j          �? H��65@�&� j        H��6E@nt� �J� j        H��6E@�l� j          �? H��65@n�� ��� b           H��65@��� b                  &ͦ ��������2       ަ ��������    Y ��   �� �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  fIDATx��?kA�ܟ����F	Wi�u���$`e%V~+?�eK!1)-m{���"j����DB����ng��͆��d�g~�����h @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @��@�Ҩ�---ݝ�������5��J��.�;������[��J��}����ˬ���i��3��) Qң}e}���s��^kķ�����g�xEHW����I�ڸ�@aX� t:����qo�j���AH�{��U�И��Z�j���}�aqq�jQ�Q��CP1 �U������6�n�_�{�Qa�:'@�X� �B���s�Hɝ�w��:��(��k�����s~������|��fى��የ������n�|�>��h�������I=��mޏi�;�t��zvb��8���Y?1����@z�^�S�UZl���cnuu�S���sL\�o�ڞ��;v�����0� �Ř��	�F��o��/
.{�� ��%m��`0����vo �Y� x� d�c7?���}R�U�P� ����&�F� Z&5@��O.�5&��q�P� T��d�Z֟��x��Ou�����x"8<x�w��ѯ42��`����Z�'�z�R�NA��h�^�m,�V��9�P忄��%��p6�JUH�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� ���ŋ8s�dҮ    IEND�B`�   g��     �� ������    R e l a t i o n a l   L i n k           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ooo�]]]�]]]�������������������������������������������������������������������������������������������������������������������������ppp�]]]�]]]�������������������������������������������������������������������������������������������������������������������������rrr�]]]�]]]�������������������������������������������������������������������������������������������������������������������������sss�]]]�]]]�������������������������������������������������������������������������������������������������������������������������uuu�]]]�]]]�������������������������������������������������������������������������������������������������������������������������vvv�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������www�]]]�]]]�������������������������������������������������������������������������������������������������������������������������yyy�]]]�]]]�������������������������������������������������������������������������������������������������������������������������zzz�]]]�]]]�������������������������������������������������������������������������������������������������������������������������{{{�]]]�]]]�������������������������������������������������������������������������������������������������������������������������|||�]]]�]]]�������������������������������������������������������������������������������������������������������������������������}}}�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�������������������������������������������������������������������������������������������������������������������������~~~�]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f�� <   �� ������ }� ��������!� ��������� Z    R e l a t i o n a l   L i n k 4   R e l a t i o n a l   L i n k [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] ~� ������ pA� �=� K    
   S�qǽr@         �|� K    -DT�!	@   
 <        ��� J   
        �?r�q_w@�̽ J           �?��8��ϐ@    �� J          �?�qǽb@�� J          �?         �q�q l@ ��8��ϐ@      _�@ ��8��ϐ@iI�          ��q��r@      �      @j~�  ���� ���� � �          �o� ������ ֿ ��������p�� ��� G   *   ��qǽr@�� O   *    X     �I@�� J    �'DT�!�? �'DT�!�? g        �/� B     Z�qǽb@�M� J     [      �9�    �s� J          �?�qǽb@��� K          �?     �9@ i�� ��� @   ~   �qǽb@�qǽb@      $@     �D@     q�      �        ��% % %                   r7�                                             sh�      A    A    A    A �       �B      �o�                       {��                           ���       |��                                       %�� ����F�  ���     �
�               ��             �����F�    r e l a t i o n a l   l i n k 9�� ������    R e l a t i o n a l   L i n k         ���     ���        <�� ������  =�� ������                       �?      �?                ?�� ������  C!� ��������                              �?        tE�          ��U U U          �?uc�   ��  ��U U U         u}�   ��    ��                                 :�� ��������                                                        ��� �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  :IDATx��1    �Om�@a��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`��0`�<0� ���b    IEND�B`�   g��     �� ����� ,   A N D   J u n c t i o n   ( p r o c e s s )           �?�   !   !                                                                                                                                       sss�\\\�^^^�^^^�^^^�]]]�]]]�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�[[[�����^^^�����������������UUU�����������������������������������������������������������������������������������������������������^^^�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������lll�[[[�___�����������������WWW�����������������������������>>>�111�SSS�������������������������������������������������������������lll�[[[�___�����������������WWW�������������������������111�kkk�����hhh�111���������������������������������������������������������lll�[[[�___�����������������WWW���������������������UUU�111�������������111�VVV�����������������������������������������������������mmm�[[[�___�����������������WWW���������������������___�111�������������111�iii�����������������������������������������������������mmm�[[[�___�����������������WWW�������������������������111�YYY�����lll�333���������������������������������������������������������mmm�[[[�___�����������������WWW�������������������������xxx�111�111�HHH�������������AAA���������������������������������������������mmm�[[[�___�����������������WWW�������������������������777�\\\�333�777���������yyy�111���������������������������������������������mmm�[[[�___�����������������WWW���������������������999�PPP���������222�999�����qqq�111���������������������������������������������mmm�[[[�___�����������������WWW���������������������111�����������������111�:::�BBB�VVV���������������������������������������������mmm�[[[�___�����������������WWW���������������������111������������������111�111�������������������������������������������������mmm�[[[�___�����������������WWW���������������������111�<<<�����������������NNN�111�===���������������������������������������������mmm�[[[�___�����������������WWW���������������������JJJ�111�AAA���������VVV�BBB�����111�???�����������������������������������������mmm�[[[�___�����������������WWW�������������������������]]]�111�111�111�[[[�������������111�BBB�������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������WWW�����������������������������������������������������������������������������������������������������mmm�[[[�___�����������������UUU�����������������������������������������������������������������������������������������������������lll�[[[�___�UUU�XXX�XXX�XXX�WWW�WWW�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�UUU�\\\�f�� 5   �� ��������b� ����b� �     A N D   J u n c t i o n   ( p r o c e s s ) ;   A N D   J u n c t i o n   ( p r o c e s s ) [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] �� ������ pv�       Y@       Y@                l@      ̐@    �K� J          �?     I@�m� J          �?      I@ i~�                 Y@�����x�      Y@ j��  ���� ���� � �          ��� ������ �� ��������p�� ��� C   *   W      @�� C   *    X   `U}I@         �A� J          �?     I@�h� B           �?   XU__@    ��� J          �?      @��� J          �?   `U}9@ i�� ��� @   ~         @      @      @   `U�G@     q!�      �        ��% % %                   rR�                                             s��     @@   @@   @@   @@ �       �B      ���      ��� ��� J                ��� J                �� ��� J            Y@�� J                �Q� �+� J                �I� J             Y@��� �l� J            Y@��� J             Y@                {��                           ���       |��                                       %� ����y�  ��     �)�               �>�             �����y�    A N D   j u n c t i o n ,   A N D   p r o c e s s 9�� ������ ,   A N D   J u n c t i o n   ( p r o c e s s )         ���     ���        <�� ������  =� �����                       �?      �?                ?-� ����-�  Cb� ��������                              �?        �� ���������� ������    f�� ;   �� ������ !� ����~� 	� ���������� ���������            � ����)� p�� �� K	            S     Y@�/� K	            S      Y@         �[� J          �?     I@�~� J          �?      I@    ��� J          �?     I@��� J          �?      I@ i�� ��� A   ~                Y@              Y@ j�  ���� ���� � �          �7� ������ j� ��������p2� �j� K            S     Y@��� K            S      Y@         ��� J          �?     I@��� J          �?      I@    �� J          �?     I@�)� J          �?      I@ iH� �F� @   ~   ������>@VUUUAQ@   @U�0@   ���T@     q��     �        ��% % %                   r��                                           & s0�  ��� B    �������?  �A�� B    �������?  �A   @@   @@ �       �B      �7�                       {v�                           �v�       |��                                       %�� ������  ���     ���               ���             �������     9� �����             ��     ��        <-� ����-�  =j� ����j�                       �?      �?                ?x� ����x�  C�� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         u	�   ��    ��                                   m~�      nt� �N� k                �l� k                n�� ��� j                ��� j             Y@n�� ��� j            Y@��� j             Y@n:� �� j            Y@�2� j                n~� �W� b                  �v� b                  &�� ��������2       f�� ;   �� ��������� ����r� �� ���������� ���������            � ������ p�� �� G    333333�?     .@�9� O	            S      Y@         �a� N                ��� N          �?      I@    ��� J                ��� J          �?      I@ i�� ��� @   ~                .@              Y@ j�  ���� ���� � �          �                     {j�                           �j�       |��                                        %�� ������  ���     ���               ���             �������     9� �����             ��     ��        <!� ����!�  =^� ����^�                       �?      �?                ?l� ����l�  C�� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                   mr�      nh� �B� k                �`� k                n�� ��� j                ��� j             Y@n�� ��� j            .@��� j             Y@n.� �� j            .@�&� j                nr� �K� b                  �j� b                  &�� ��������2       �� ��������       ���   ��� N  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�]�K��'�0'�LgTEPΜs(�1��Cŀ"�3�z&�s�{��̟�{v��9��]�lO�z��]]]K�Hq@q@q �̂v��-���Os\�ᧁr#,�������hbb�K4�^o/!!a] < >>>E�������Qqqq����#�B�KC|��=*99?��h� A ��Y�f)�����)\�޽;6,6&&&ܢ*�_�@RR-^����T:=�������7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ���7F�@`�Bހ�g�/���F>|�w��Q�c*T�bcc}9�H�;���ХK�����t���w�fʑ#+V��-J�K��6m�P����Y�
���c�h�ƍt���߿O�\�~]˷e��۷/u�Ё2f��-��D_�	0�\��رc`'�O�>�ҥK��СCvY|'�L���+�ի=�<ՂB'N$�	_����3^ӦMs@���T�RT�D	J��y�˖-����˂� ���z�Νp���w޼y5�ԬY�2dȠ�����۷�V�XA_�~e�]�hիW�r�����矅GGz��}Z�|9�w5j� ��nݺ �9S�LԾ}{ڽ{�63�*���#m۶���xaA�n�:���02g�L�g����,H3g���=j[��"���o��ԩSLY��ٓ����L�*U��m�g��ӧO��K��5�W�B� ����v� Z�l�L�&ԩS�􌝂�IH�e��P�dɒܬ�A�����7o�r�k �m�^v<�A�,$��c��ϟYI��<@�@8��mD
	�`p&��{�@��'OĘ�.
	�
pG�k�.n�9'�,*_�<EE��߀X�{&^H.\�+�;vЗ/_�����:u��L�S�� �QH�&M�r�+aܸq���of$9r�y�?~jڴ)��_��ߥK�0�ϙ3����ݻ�Ɛ��k׮��'HXT�V�p>�#�3�`/`�/^ШQ��G;jѢu���.ɗq Ҙ?>a}�#Xu�ؑnܸA�>�Z�J3y��m�F�ь3�kۂG
=��G�8+����2��H�=�Q��Z�ji��{ܺu�Ν;g[��V�Z٦�)4�`�l޼�F�M�?����0@�&� *�z��8���B�t��bx���T�~}=*�o�����{��.���+	?肁R'\=��y�q��z�~�b&�|��fp����9y�dm�J!��s�p��������w�҇�h�2�n޼�˦��@�-[6��^� 4`����Z�hƢ<`�8x�`JNN�e�j��K�D\�>}�- bbbhӦM��Võk��v���"������n��3��x��M�X Ν;�ʔ)��; �.r�.������ѣG�8���w�m[��"��ʕ+m �v�֍6l�f��<�jժA�����ߟ``j%ީ$t"�p ���g����� �eɒ� �ʕ+�%q02���޾}k��I�g�E�[��ܹs��)k֬��AŊ�y�  @�h�:z���m���h*^��m�(�B���������`�Eܚ5k�\�rA��0��[�afѯ�Y�Dy
�{���;���B�fq�ڵ��
=����Ç�hd� >>ޮ�PqB� �)R�������\esz�cۈ��,+f+g��ٺX37�{9W�\�~�z�u��.k��m���ֺ��,�L �A��"�� � 6l �$����`� ��9���"͉pk	3B8J>��@ [1|X���[2+�5 �� +�PG��&�:��#��;�E���[3�ʙ�a����~"�`���L�z�`$r<��&�3���!vNm�d}����+��z�
p>ɣիWk�	yyBIöq���Y�e��:�c�c� ��G8橕ye�iP��1�2�6�e��$B1$ݻw/]�r%by@)4bĈ��'O��	&pO"��_((��ECK!\J��8���ڵkڶ/))���6����4e���m!�D
��R����U�p�B�Z(�S�U�ޠO�>�3 v%�f�"X,�����Lk'^9�ӄ39/[�,AS�{�Nt��j۶�fC�r�� Ϧ8l�11�GN�8A/^d�8~Ƃ�B�
�^`�С��a�0i�$G�:��o�0��q����N��<��O�a��-  �^�:-Y�D��x�={�h@��mH����s�i˘`��+%...����EX�u5=3������˸�-$�,\Fݺu+9�!���U�T�\�6h���8T���tx��0`�:	0@�Us��c�N-A��&�W�S��͛�ԩS���;����$4�X7��{�Q ��p	�ɸ���� ��\7��ha�t��msQO��\�q�#G�Ԅe��NQ���npaZ��B|p
�t�RB��mxL�Gd�t!`&�z٪b�~�#\FQ�߁ xx�=�k��j�WH�5�����h�ủZU �8���;|�T�
��;�Q p��jU��S�p�3
���S�*xJ�tF���{�UO�Ý�(��wO��@�)q��w��V<%w:�@��=ժ����Ng�ủZU �8���;|�T�
��;�Q p��jU��S�p�3
���S�*xJ�tF���{�UO�Ý�(��wO��@�)q�ә�[�Ϟ=K��x}pK����?�z�w�p .���	 Jo&��I������w�O+�<�����*��x^��qXp�33m[R�+(�Á��\0�%��    IEND�B`�   g�#     �# �����# *   O R   J u n c t i o n   ( p r o c e s s )           �?�   !   !                                                                                                                                       ]]]�^^^�^^^�^^^�\\\�\\\�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�]]]�___�����VVV�������������������������������������������������������������������������������������������������������������������������bbb�]]]�```�������������������������������������������������������������������������������������������������������������������������ddd�]]]�```�������������������������������������������������������������������������������������������������������������������������ddd�]]]�```�������������������������������������������������������������������������������������������������������������������������ddd�]]]�```�������������������������������������������������������������������������������������������������������������������������eee�]]]�```�������������������������������������������������������������������������������������������������������������������������eee�]]]�```�������������������������������������������������������������������������������������������������������������������������eee�]]]�```�������������������������������������������������������������������������������������������������������������������������fff�]]]�```�������������������������������������������������������������������������������������������������������������������������fff�]]]�```�������������������������������������������������������������������������������������������������������������������������fff�]]]�```�������������������������������������������������nnn�DDD�111�:::�aaa�����������������������������������������������������ggg�]]]�```���������������������������������������������888�111�XXX�}}}�eee�666�111�������������������������������������������������ggg�]]]�```�����������������������������������������===�333���������������������FFF�111���������������������������������������������ggg�]]]�```�����������������������������������������111�{{{�������������������������111�TTT�����������������������������������������ggg�]]]�```�������������������������������������bbb�111�����������������������������DDD�111�����������������������������������������hhh�]]]�```�������������������������������������EEE�111�����������������������������ccc�111�����������������������������������������hhh�]]]�```�������������������������������������111�999�����������������������������uuu�111�����������������������������������������hhh�]]]�```�������������������������������������???�111�����������������������������ggg�111�����������������������������������������hhh�]]]�```�������������������������������������\\\�111�����������������������������KKK�111�����������������������������������������hhh�]]]�```�����������������������������������������111�����������������������������111�HHH�����������������������������������������iii�]]]�```�����������������������������������������666�777���������������������SSS�111���������������������������������������������iii�]]]�```���������������������������������������������111�222�vvv���������BBB�111�fff���������������������������������������������iii�]]]�```�������������������������������������������������LLL�111�111�111�===�����������������������������������������������������iii�]]]�```�������������������������������������������������������������������������������������������������������������������������jjj�]]]�```�������������������������������������������������������������������������������������������������������������������������jjj�]]]�```�������������������������������������������������������������������������������������������������������������������������jjj�]]]�```�������������������������������������������������������������������������������������������������������������������������jjj�]]]�```�������������������������������������������������������������������������������������������������������������������������kkk�]]]�```�������������������������������������������������������������������������������������������������������������������������kkk�]]]�]]]�������������������������������������������������������������������������������������������������������������������������kkk�]]]�UUU�XXX�XXX�XXX�UUU�WWW�XXX�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�UUU�sss�]]]�f� 5   � ��������� ����� 4     O R   J u n c t i o n   ( p r o c e s s ) :   O R   J u n c t i o n   ( p r o c e s s ) [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] � ���� p�       Y@       Y@               �u@      ̐@    �� J          �?     I@�� J          �?      I@ i�         @_�     Y@�����x�      Y@ j�  ���� ���� � �          ��	 ����@ 3	 ��������p� �7 C   *   W      @�X C   *    X   `U}I@         �� J          �?     I@�� B           �?   XU__@    �� J          �?      @�� J          �?   `U}9@ i	 �	 @   ~         @      @      @   `U�G@     qc	      �        ��% % %                   r�	                                             s�	     @@   @@   @@   @@ �       �B      ��	      �
 ��	 J                �	
 J                �R
 �,
 J                �J
 J             Y@��
 �m
 J            Y@��
 J                ��
 ��
 J            Y@��
 J             Y@                {                           �       |@                                       %N �����  �W     �k               ��             ������    O R   j u n c t i o n ,   O R   p r o c e s s 9 ���� *   O R   J u n c t i o n   ( p r o c e s s )         �     �        < ����  =[ ����[                       �?      �?                ?i ����i  C� ��������                              �?        � ��������� �����    f� ;   � ����� ] ����� E ��������� ��������5            W ����e p �? K	            S     Y@�k K	            S      Y@         �� J          �?     I@�� J          �?      I@    �� J          �?     I@� J          �?      I@ i" �  A   ~                Y@              Y@ jW  ���� ���� � �          �s ����� � ��������pn �� K            S     Y@�� K            S      Y@         �� J          �?     I@� J          �?      I@    �C J          �?     I@�e J          �?      I@ i� �� @   ~      @>@   �}Q@   @U�0@   ���T@     q�     �        ��% % %                   r                                           O sl  �/ B    �������?  �A�M B    �������?  �A   @@   @@ �       �B      �s                       {�                           ��       |�                                       %� ����,  ��     �               �#             �����,     9[ ����[             �N     �[        <i ����i  =� �����                       �?      �?                ?� �����  C� ��������                              �?        t          ��U U U          �?u+   ��  ��� � �         uE   ��    ��                                   m�      n� �� k                �� k                n� �� j                �� j             Y@n4 � j            Y@�, j             Y@nv �P j            Y@�n j                n� �� b                  �� b                  &� ��������2       f� ;   � ��������Q ����� 9 ��������� ��������6            Y ����� p �I G    333333�?     .@�u O	            S      Y@         �� N                �� N          �?      I@    �� J                � J          �?      I@ i$ �" @   ~                .@              Y@ jY  ���� ���� � �          �                     {�                           ��       |�                                        %� ����   ��     �               �             �����      9O ����O             �B     �O        <] ����]  =� �����                       �?      �?                ?� �����  C� ��������                              �?        t          ��U U U          �?u   ��  ��� � �         u9   ��    ��                                   m�      n� �~ k                �� k                n� �� j                �� j             Y@n( � j            .@�  j             Y@nj �D j            .@�b j                n� �� b                  �� b                  &� ��������2       � ��������       ��   ��# �
  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  
IDATx�]g���5�(��PQT�9�YWT"�
��#�̫�	T�����pq��s\��7ܖsu���	�ӧ��лS���s��A )�>}�,�����,�����:�<�$����9rJMM}��r�,�w�7�Y�f�Y���ӧ��4i���(�$$^���K�۷o��d�d�Ju��9#%%�_�e�%''ӄ	
�ɓ'�Q%�\�z��-[�Ue%��B�b_H`��UՅ
	�}!���WU($,��+_U]H����X�|Uu!�B�b_H`��UՅ
	�}!���WU($,��+_U]H����X�|Uu!�B�b_H`��UՅ
	�}!���WU($,��+_U]H����X�|Uu!�B�b_H`��UՅ
	�}!���WU($,��+_U]H����X�|Uu!�B�b_H`��UՅ
	��_6�l��������Kz��,X�J�,I�
���V���͛t��1r��ѳg�\�;��Px޼y�D�T�tijР�iӆ�֭K�n�-aIp��}ںu+?~�U����ׯ_�ɓ'����˴q�F*^�8�jՊz��E����$����o޼�իW�Ν;)===j�~�������:t�@�Ǐ�
*D�n�H���cA�6m�D=z���۷Ǆ �+����ԻwoZ�|9��H�$�?o�<h�>�U7߾}�6И1c����q�˯č'��I�&Ѿ}���������4|�pz�Ⅿ��#3���;���p]ժU�e˖T�|ywZX�H��铫L�N�:Eׯ_+9�>0:�֭[G�ʕ+NM�+V�E �X<x0u�҅@΁T�?&��h�uM>�Κ5�֮]K�}h.��ʌ�Ν;G�7o�۸qcڱc�ۇ����o��ݻ]��^>Z"JMuF� ��ܹs��4�֬YCU�Tц�, �.\H,о�h��ݻ�Y2�f$	V�\�6�������'rAu�ڕfϞ͆Ǭa���l��
�#�h4Ӝk߾=M�2��eVǍ���*�+W�0AG��{�6�6��N��m���sχBիW炸Ul� 
�"�ϟ?�A�#F�����r��I3f�`�Ƭ�իWl��	�"��'(--��ʕ+��-'Oy,�Dj۶�gR?~��]�vyʃ(0�G�a1�޽�/۾؟��ѣG9q�dF��ҥK,�X��5oޜ�rp~���QƬ�a	pg�\Æ}��͕+9_��*���y��5Oy�Ɛ �/�5mڔ�\�|��MS�j��}C�5k���Z�j�����F�Yh	�޽�B�S
9a�2e�q��;w"H5{�C�	��B)~;�x\y�.�.?cH�m�V�TIWϸ�+V���Ǐ�r��3�(Ɛ�{��뾀._��Q�,�Q�Q@�#G�(��yT#H��Xn�7����H -A���m��������o�N6s����addDK�?~�*���*P� [�� �p9�1���'�MpF� @r��/E����*S$�C�{�O�ψQ
t���Qf��Ɛ�{�<x3@���/`ʕvcHP�X1O��}���>}�)�� ����MqƐ�[��7n��s\Y�5x/W�vm/Q��C�z���qo%1B�.?]y#�6.ь!A�:u�>I�t���q���3�8���50�6:t�g-q��C.��	C`LK���l�e� ����!��s��`1�;vdQۿ?���F΂055��Be#f��(���%�.�U��
%���g�z��\`5�E ��Ɯ۲eݺu��[�K�.e�w�֍��`#g��8���ca�jΜ9l�	ְ��h�"���~��E�|��1��%0�-.�E, cd�kݺ5U�V�D�q$ �#F�`���*�'���!��}���mt6�-J3g��%H��$��&dp�s.\p�Ob���x�"8е����*UJ,�r#I $kԨA�G�ւ�� c��:����|Þ>}:6,�(�ڵk�-KP�RPK�O�`9��Ж��C�ѨQ#�-��h�1vx���k�̙3YT"�iӦi�r �I�cg0���h���e���/ZS��/&,����0 9y�d5j�z�߳gOZ�d�� XF���9r�;N�����b�7�`,o�81-�&��!��E��m�6��,�ɣ��1�����L)))ƭ�Q��$	P7La���`�#}�
����Al|�lٲ����&	�Zp&��p'��ɓ�`� l4���j��"�"<Lߩo �&2ZS��
�p��%Ah�1{�ԩ��}��`�^�56SN��?V[A/�0�0媘Wb���)b,@�=!��p�/$	���; ��i	�����	�Bဴ���@@��!�p@Z�t�  cၐ@8 -�p@�� �1��@H ��@8 ݁p Ș@x $HK p�׭�G��q�pÝ���4�̽�[�D��g�T�����_��������Y��s�?ݹ��,��/�8��8���~��E��IRs�7���c�    IEND�B`�   gY     Y ����Y 0   S y n c h r o n o u s   A N D   J u n c t i o n           �?�   !   !                                                                                                                                       rrr�\\\�^^^�^^^�^^^�]]]�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�\\\�VVV�^^^�^^^�^^^�[[[�����^^^�����������������UUU�����������������������������������������������������������������������������������������������������]]]�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������>>>�111�SSS�������������������������������������������������������������kkk�YYY�___�����������������UUU�������������������������111�kkk�����hhh�111���������������������������������������������������������kkk�YYY�___�����������������UUU���������������������UUU�111�������������111�VVV�����������������������������������������������������kkk�YYY�___�����������������UUU���������������������___�111�������������111�iii�����������������������������������������������������kkk�YYY�___�����������������UUU�������������������������111�YYY�����lll�333���������������������������������������������������������kkk�YYY�___�����������������UUU�������������������������xxx�111�111�HHH�������������AAA���������������������������������������������kkk�YYY�___�����������������UUU�������������������������777�\\\�333�777���������yyy�111���������������������������������������������kkk�YYY�___�����������������UUU���������������������999�PPP���������222�999�����qqq�111���������������������������������������������kkk�YYY�___�����������������UUU���������������������111�����������������111�:::�BBB�VVV���������������������������������������������kkk�YYY�___�����������������UUU���������������������111������������������111�111�������������������������������������������������kkk�YYY�___�����������������UUU���������������������111�<<<�����������������NNN�111�===���������������������������������������������kkk�YYY�___�����������������UUU���������������������JJJ�111�AAA���������VVV�BBB�����111�???�����������������������������������������kkk�YYY�___�����������������UUU�������������������������]]]�111�111�111�[[[�������������111�BBB�������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������kkk�YYY�___�����������������UUU�����������������������������������������������������������������������������������������������������jjj�YYY�___�UUU�XXX�XXX�XXX�WWW�XXX�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�XXX�UUU�XXX�XXX�XXX�UUU�[[[�f�L 5   �L ��������V; ����V; �     S y n c h r o n o u s   A N D   J u n c t i o n =   S y n c h r o n o u s   A N D   J u n c t i o n [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] �6 �����6 ph6       Y@       Y@               �}@      ̐@    �=6 J          �?     I@�_6 J          �?      I@ ip6         @o�     Y@�����x�      Y@ j�6  ���� ���� � �          �|8 �����9 �7 ��������p�7 ��6 C   *   W      @�7 C   *    X   `U}I@         �37 J          �?     I@�Z7 B           �?   XU__@    ��7 J          �?      @��7 J          �?   `U}9@ i�7 ��7 @   ~         @      @      @   `U�G@     q8      �        ��% % %                   rD8                                             su8     @@   @@   @@   @@ �       �B      �|8      ��8 ��8 J                ��8 J             Y@�9 ��8 J                ��8 J                �C9 �9 J            Y@�;9 J                ��9 �^9 J            Y@�|9 J             Y@                {�9                           ��9       |�9                                       %�9 ����i:  �:     �:               �0:             �����i:    s y n c h r o n o u s   A N D   j u n c t i o n 9�: �����: 0   S y n c h r o n o u s   A N D   J u n c t i o n         ��:     ��:        <�: �����:  =; ����;                       �?      �?                ?!; ����!;  CV; ��������                              �?        �L ��������oL ����oL    f�B ;   �B �����B A ����rB �@ ���������@ ���������            = ����= p�< ��; K	            S     Y@�#< K	            S      Y@         �O< J          �?     I@�r< J          �?      I@    ��< J          �?     I@��< J          �?      I@ i�< ��< A   ~                Y@              Y@ j=  ���� ���� � �          �+? �����? ^> ��������p&> �^= K            S     Y@��= K            S      Y@         ��= J          �?     I@��= J          �?      I@    ��= J          �?     I@�> J          �?      I@ i<> �:> @   ~   ������>@VUUUAQ@   @U�0@   ���T@     q�>     �        ��% % %                   r�>                                           & s$?  ��> B    �������?  �A�? B    �������?  �A   @@   @@ �       �B      �+?                       {j?                           �j?       |�?                                       %�? �����?  ��?     ��?               ��?             ������?     9@ ����@             �@     �@        <!@ ����!@  =^@ ����^@                       �?      �?                ?l@ ����l@  C�@ ��������                              �?        t�@          ��U U U          �?u�@   ��  ��� � �         u�@   ��    ��                                   mrB      nhA �BA k                �`A k                n�A ��A j                ��A j             Y@n�A ��A j            Y@��A j             Y@n.B �B j            Y@�&B j                nrB �KB b                  �jB b                  &�B ��������2       f{G ;   {G �����G 	F ����fG �E ���������E ���������            D �����D p�C �C G    333333�?     .@�-C O	            S      Y@         �UC N                �xC N          �?      I@    ��C J                ��C J          �?      I@ i�C ��C @   ~                .@              Y@ jD  ���� ���� � �          �                     {^D                           �^D       |�D                                        %�D �����D  ��D     ��D               ��D             ������D     9E ����E             ��D     �E        <E ����E  =RE ����RE                       �?      �?                ?`E ����`E  C�E ��������                              �?        t�E          ��U U U          �?u�E   ��  ��� � �         u�E   ��    ��                                   mfG      n\F �6F k                �TF k                n�F �xF j                ��F j             Y@n�F ��F j            .@��F j             Y@n"G ��F j            .@�G j                nfG �?G b                  �^G b                  &{G ��������2       foL ;   oL ���������J ����ZL �J ���������J ���������            I �����I p�H ��G G    333333�?     .@�!H O	            S      Y@         �IH N            Y@�lH N          �?      I@    ��H J            .@��H J          �?      I@ i�H ��H @   ~                .@              Y@ jI  ���� ���� � �          �                     {RI                           �RI       |�I                                        %�I �����I  ��I     ��I               ��I             ������I     9�I �����I             ��I     ��I        <	J ����	J  =FJ ����FJ                       �?      �?                ?TJ ����TJ  C�J ��������                              �?        t�J          ��U U U          �?u�J   ��  ��� � �         u�J   ��    ��                                   mZL      nPK �*K k                �HK k                n�K �lK j                ��K j             Y@n�K ��K j            .@��K j             Y@nL ��K j            .@�L j                nZL �3L b                  �RL b                  &oL ��������2       �L ��������       ��L   �Y s  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�]���>k�����)�^AQ|*����(v�^�`��
���>�`Wt-�6�X֮����#�s�g&��}��d��%���s�;�r�	�"��Ł+���$''���E���y���(����Oc5����#��_�~-NHH��i�b ��5Эv���F\�׳g��ԬY3I�/�*T9ܼy3S�b�ReȐ�!5��/_�Н;w�i%����@���Ϳ4���ڷo�����ף*�@|||�k�B#��KLLL�իW��TF@]�����7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ���7{�@`�Bހ�*�,мt������۷���*P� e͚5�ݍ�_���ǉ.\�@'O��S�Nѽ{�@�R�l٨H�"T�pa*Y�$�iӆbcc�Y�
��#Ghݺup���w��+W���6n�H}��!���K��[6����`�:t(�3� NBLJJ�E��#��:N����˗ԳgOz��Y��:&L�@��[7�z���	�
�2e�+ ҤIC%J� �(�J���ŋ�޽{�@��K�G��۷��B�)�ܹs� �Q��M�?��߾}�ݻw�ҥK����̲,�z��Q��ٙy������iO�߿OK�,a>]���	 �[��	 dN�>=�k׎v�ܩ��
>|�@[�la%*^X�^�����(8��9s&�_�?~�>}:��p��a���)$��ĉLY��у����L7*T��/�{���ӧ���{t����_�~e
�E��4{����r��B�IH�����R��ŹY�t�_�f���p��FXA�H��d!A����Ǐy2�[P�ɨ���<��L �!��j��B�\�e�)$������;���D�4��lٲ$�w��A����ٶm}��%[3�����3�큎;ڣy/$�ҤI�@�J;v,i�b�A¡C���y�楦M�r�%QH���;w�� ���Y��y�޽���2t�҅p�$	�*U��x���ѣG�����s9r$a�щ�7oN�:urJ
d�� �4�ΝK���F:t��W���˗/וG�<y�X�Q�F4m�4�ñ���B�w8�ő0�
��v�L�,ҽ{wk�cX���,�׀�uR:s�c9,#[�l�&B��  ��(�a�5j=~�8*�c?����6� P�K�t�95���� �u`�[�n����Qa]�[ Mc�h���N��*	?���N���s�̡ƍUH{�Hp��E]/`���	rҤI��1�Bv�k�H����{�졾}�27}x��������ƍ�lzY��~�޵2�e��r��}�]�y���ʢ<�c�8h� �}�6/w�Q��˺ߗ#��S�: S�L�~�z}�Zõj��>NHP^eoZt�F!G���>w�1A�={6�*UJ�'V �.r�]����ѣG�8���w��X��"���e� �v�ڕ6l�f(�@=�r��!��(���׏�`j'ީ$�*D&�@ ��ӧO;��� �e̘� ��+:%�qP2�fmo޼1��
v���{�E�Z���9s��)s����A���y�  `Ѫu���+�2�S���E�:��)�H�� Ü܉�qqqN�!q�ĭ\��ʔ)o���`� �՞#�a�fO�^(�����>n;��V��TqNׇ�@����:u�8*N(`>��B�
q������ln�s,a���bV �s�7��'k��y/�ȑ�֬Y�����e��� ����^��	�;�"�-���v�Z�H)a"*���,�Y�RCGX�V����0"D�����QH`)��<xฅ��o� 0"@�8�t$�	�N��l��"X)���r�x�+bDp�OD�<���Z��� ��D�G<k"^9k�b���Tև�5�����P ��I�X�B�O��N���ƍs͊%+T�YS\+�I�@ �C<0o[�W֚��!�<�C�@�m\�JB� E҄�JLL�Z�>|xD��Ǐ���㹊'Q?�?PP(`)�4�`��q����˗�e����y�ӎ=J����#n�B>�
���n���U8�|][(�SXU@ߠw�ގ# V%3f� h,�����Lm'^9�ӄS9/]�4a�v�nt��9j۶��C�r�O�gS6��#ǎ����3G?c�Y�\9}_`Ȑ!����0q�DW��=�?�.����`��n��<��_�a��-  �Z�*-\�P�x�]�v�@��mH����s�mɘ`��+�Z�j!���aY�jFfxSw�a���*$�,�nڴ���F��J�*�.q4h�X[���vx��P`�;	0@��9��1t�� Th����T�Y�f4y�d�&���q�����	����(�FJ8N��:S�A��nLP��Y�ӭ[��E}rb��A(��1B"6�0�99D�f���jN
��) ���J	W����1?�)0 0��� ���-f��c��(�B98�vﯻ�ǜ�ڂ~N,qx�o��V|%oF�����U_�Û�Q ���jU��W���a�ữZU �8�yo��V|%oF�����U_�Û�Q ���jU��W���a�ữZU �8�yo��V|%oF�����U_�Û�Q ���jU��W���a�ữZU �8�yo��V|%oF�����U_�Û�	�J�wR�2���W�z���7�Q�P��&��TF��J1�M�֭�i��4��?��\Qǋ�WE8���b��>dq���P4$J�ՐZs��_�-ϿCԍ����"G��M�    IEND�B`�   gߌ     ی ����� .   S y n c h r o n o u s   O R   J u n c t i o n           �?�   !   !                                                                                                                                       ]]]�^^^�^^^�^^^�UUU�\\\�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�___�^^^�^^^�^^^�]]]�```�����VVV�����������������������������������������������������������������������������������������������������UUU�����������������```�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������bbb�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ccc�]]]�aaa�������������������������������������������������nnn�DDD�111�:::�aaa���������������������������������^^^�����������������ccc�]]]�aaa���������������������������������������������888�111�XXX�}}}�eee�666�111�����������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������===�333���������������������FFF�111�������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������111�{{{�������������������������111�TTT���������������������^^^�����������������ccc�]]]�aaa�������������������������������������bbb�111�����������������������������DDD�111���������������������^^^�����������������ccc�]]]�aaa�������������������������������������EEE�111�����������������������������ccc�111���������������������^^^�����������������ccc�]]]�aaa�������������������������������������111�999�����������������������������uuu�111���������������������^^^�����������������ccc�]]]�aaa�������������������������������������???�111�����������������������������ggg�111���������������������^^^�����������������ccc�]]]�aaa�������������������������������������\\\�111�����������������������������KKK�111���������������������^^^�����������������ccc�]]]�aaa�����������������������������������������111�����������������������������111�HHH���������������������^^^�����������������ccc�]]]�aaa�����������������������������������������666�777���������������������SSS�111�������������������������^^^�����������������ccc�]]]�aaa���������������������������������������������111�222�vvv���������BBB�111�fff�������������������������^^^�����������������ccc�]]]�aaa�������������������������������������������������LLL�111�111�111�===���������������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ccc�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ddd�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ddd�]]]�aaa�����������������������������������������������������������������������������������������������������^^^�����������������ddd�]]]�^^^�����������������������������������������������������������������������������������������������������ZZZ�����������������ccc�]]]�UUU�XXX�XXX�XXX�UUU�WWW�XXX�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�ZZZ�WWW�XXX�XXX�UUU�jjj�]]]�f� 5   � ���������p �����p      S y n c h r o n o u s   O R   J u n c t i o n <   S y n c h r o n o u s   O R   J u n c t i o n [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] l ����l p�k       Y@       Y@               ��@      ̐@    ��k J          �?     I@��k J          �?      I@ i�k         pw�     Y@�����x�      Y@ jl  ���� ���� � �          ��m ����Yo Lm ��������pm �Pl C   *   W      @�ql C   *    X   `U}I@         ��l J          �?     I@��l B           �?   XU__@    ��l J          �?      @�m J          �?   `U}9@ i*m �(m @   ~         @      @      @   `U�G@     q|m      �        ��% % %                   r�m                                             s�m     @@   @@   @@   @@ �       �B      ��m      �*n �n J                �"n J             Y@�kn �En J                �cn J                ��n ��n J            Y@��n J                ��n ��n J            Y@��n J             Y@                {(o                           �(o       |Yo                                       %go �����o  �po     ��o               ��o             ������o    s y n c h r o n o u s   O R   j u n c t i o n 9-p ����-p .   S y n c h r o n o u s   O R   J u n c t i o n         � p     �-p        <;p ����;p  =xp ����xp                       �?      �?                ?�p �����p  C�p ��������                              �?        � ��������ԁ ����ԁ    f�w ;   �w �����w zv �����w bv ��������v ��������            tr �����r p(r �\q K	            S     Y@��q K	            S      Y@         ��q J          �?     I@��q J          �?      I@    ��q J          �?     I@�r J          �?      I@ i?r �=r A   ~                Y@              Y@ jtr  ���� ���� � �          ��t ���� u �s ��������p�s ��r K            S     Y@��r K            S      Y@         �s J          �?     I@�:s J          �?      I@    �`s J          �?     I@��s J          �?      I@ i�s ��s @   ~      @>@   �}Q@   @U�0@   ���T@     q�s     �        ��% % %                   r$t                                           O s�t  �Lt B    �������?  �A�jt B    �������?  �A   @@   @@ �       �B      ��t                       {�t                           ��t       | u                                       %u ����Iu  �u     �+u               �@u             �����Iu     9xu ����xu             �ku     �xu        <�u �����u  =�u �����u                       �?      �?                ?�u �����u  Cv ��������                              �?        t*v          ��U U U          �?uHv   ��  ��� � �         ubv   ��    ��                                   m�w      n�v ��v k                ��v k                nw ��v j                �w j             Y@nQw �+w j            Y@�Iw j             Y@n�w �mw j            Y@��w j                n�w ��w b                  ��w b                  &�w ��������2       f�| ;   �| �����| n{ �����| V{ ���������z ��������            vy �����y p*y �fx G    333333�?     .@��x O	            S      Y@         ��x N                ��x N          �?      I@    ��x J                �!y J          �?      I@ iAy �?y @   ~                .@              Y@ jvy  ���� ���� � �          �                     {�y                           ��y       |�y                                        %z ����=z  �z     �z               �4z             �����=z     9lz ����lz             �_z     �lz        <zz ����zz  =�z �����z                       �?      �?                ?�z �����z  C�z ��������                              �?        t{          ��U U U          �?u<{   ��  ��� � �         uV{   ��    ��                                   m�|      n�{ ��{ k                ��{ k                n| ��{ j                ��{ j             Y@nE| �| j            .@�=| j             Y@n�| �a| j            .@�| j                n�| ��| b                  ��| b                  &�| ��������2       fԁ ;   ԁ ��������b� ������ J� ��������� ��������            j~ �����~ p~ �Z} G    333333�?     .@��} O	            S      Y@         ��} N            Y@��} N          �?      I@    ��} J            .@�~ J          �?      I@ i5~ �3~ @   ~                .@              Y@ jj~  ���� ���� � �          �                     {�~                           ��~       |�~                                        %�~ ����1  ��~     �               �(             �����1     9` ����`             �S     �`        <n ����n  =� �����                       �?      �?                ?� �����  C� ��������                              �?        t�          ��U U U          �?u0�   ��  ��� � �         uJ�   ��    ��                                   m��      n�� ��� k                ��� k                n�� �р j                �� j             Y@n9� �� j            .@�1� j             Y@n{� �U� j            .@�s� j                n�� ��� b                  ��� b                  &ԁ ��������2       � ��������       ��   �ی �
  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  
KIDATx�]g�K�3�g�
�Q1+�
�,bĀ*�ᇘ3*(��O1�`�	��CTT�3�9�'�gΞ��|���۩���ݝZ�a�ݩ����]C�IP�� �3'''O������(�EC#���Z���ݻ�~�T>�p�=%%eH�V�r�H�ϝ;�ҢE�����r��~�zj͚5S
,:C�G?}�Dw���d�~����}����'�*���3���-�9s��ܺu+�0G333s������>���OD@I �h���$���@}J�F�]e%�mD�S4��*+	l#*P��@��lWYI`Q����f��Jۈ
ԧ$h4�UV�FT�>%�@�ٮ���6��)	�v����OI �h���$���@}J�F�]e%�mD�S4��*+	l#*P��@��lWYI`Q����f��Jۈ
ԧ$h4�UV�FT�>%�@�ٮ���6��)	�v����OI �h���$���@}n�*����ʟ?��/_һw�(55�J�.ME��J���IO'��<y���j���3��_�|����T�RT�lYjܸ1u�Ё4h@y�$��LJ<x���hlt��)����x��������s��Uڼy3�,Y�ڵkG����F��(����o޼����Ӟ={�ǏQ[���״�~�ӥK�2e
U�T)j�~S���	�G[�l�>}��Ν;��wC;v����O�W�&x�dJ�I�;~ѢE�j�*���CLm���WڴiM�8�޿O����I�;rڴit�����w�/^�1c�Ћ/~��/�O���I�	7U�^�ڶmK+Vt��ŋ'���11r8{�,ݸq#,uw�ܡQ�FQFFU�P!�2~�$�k֬	� 
�#FP�=$�H���cB��or��;o�<ڸq#9�9վ��l.\�@[�n5۬Y3ڵk�ۆ�P��?��}����	���'B�TrG��1>|8mذ��U�f�*&��.]JK�,1���J������P�|}L	֮]�l����ԩS�,a�z��I���g�c԰x�b6����H�6n�K�;w�3fpYr-Ì��ɓ�r�e�v��ǯBQ$8p� ��W�C��3gݷWy��ȑ#�V�Z\w����S�8oUq;y��ݣ-�Eʛ7/9oaUcT���+6��bHp��i����İjժx���܆ �:v�������`�S�W�?~�Űw��qy��\:q�'��L	�\���ɠx�֭[�M�/p��x�1��A� ��ԤI��=�͗/u��ݫ*�L��u�r?
D� �/.�lْ[�5oޜ�i�Zl�E��j�:u�
]ݺu����N�P	�ݻ�Bc2
[8a�r��~����&���O���F�w���7���|"H�=ҭR�J8�i=O�ʕ=u~��1&K�<O�@	�;+Q�L���ͬWD��q#<e̊�����&_��(�D��j�P��B�
���o��f��q�d�'�'(\�0{)��䁊)���OBߓ �p9��OD2�+��$ߓ @r���+C���α�S�zE��X�b��g2�g�(��:�Q��jq$�Z$\e�yA I[�E��D���y��-=}��S+�x%LeKJ"H����7o�slY�6x�T�^=/�/�� AÆY𸻒-��t>S}#<m̊� A����6I�L�S���0���c9W���a��ѣG=�`��ų2a
Dx\�)fP�b`517<D ��a��lbHеkW�C����¹�޽���-Be&P(�+�5	�K�nݺ�B�f 33��x^��Ғ X�6�Ҷm�����\��ex4�r�J�|�^���l�
E� ����E��mv$X#:ڲeˌ1�����E��O���fa#� Vq��V]���F�l�
E�  �;�� 6� � 7��|����7��b"����ܹsM�|+G�B���t��%7�$F��˗/�СC�訦� @�2eL�|+G Y�vm�0a�Tx�s��u��{��ٔ���F�:u2�������5G��>|�XKD�ޣiӦ�X�s���wx���������TB׬Y����{�$��3��ZD4'a�2B��mB(��˗���'��A t��>}:�?>p(.�}���+V$ �XOl�q�ƹ��~��Q���o,A_$�aq�V:eIA\'�s�6mhǎn�Y�!O��'ފ2l�0=z����\L�?IC\���c��Ew��>bD�<D@l��|��!�K�CIE��I�&�|�'�̙3ng� <hB�9��E,E~���	1��U$��X��$�p��u��~��c:����M����k��;�I�F���y]��㢇�6 PDJe��@9��@9� �́�@I�PO���@9 �O�<P(�(�9P �(����m�@@��%�r@=�r@�� �>��@I�PO���@9 �O�<P(�(�9P �(~�����"��N��ʖ�ܜ3��"�
�-�����l�O	����������?섍�,���w�����b8��Ҝ���RMr^ڑ�y��ތ�����Ѳ��"�l���5����    IEND�B`�   gۺ     ׺ �����    X O R   J u n c t i o n           �?�   !   !                                                                                                                                       qqq�\\\�^^^�^^^�^^^�]]]�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�^^^�\\\�����___�����������������UUU�����������������������������������������������������������������������������������������������������\\\�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�```�����������������UUU���������������������~~~�QQQ�������������������������RRR�___�����������������������������������������jjj�[[[�```�����������������UUU�������������������������111�===�����������������ggg�111���������������������������������������������jjj�[[[�```�����������������UUU�����������������������������111�|||�������������111�ccc���������������������������������������������jjj�[[[�```�����������������UUU�����������������������������BBB�111���������CCC�666�������������������������������������������������jjj�[[[�```�����������������UUU���������������������������������111�TTT�����111�����������������������������������������������������jjj�[[[�```�����������������UUU���������������������������������eee�111�111�SSS�����������������������������������������������������jjj�[[[�```�����������������UUU�������������������������������������111�111���������������������������������������������������������jjj�[[[�```�����������������UUU���������������������������������ttt�111�111�TTT�����������������������������������������������������jjj�[[[�```�����������������UUU���������������������������������111�```�ddd�111�����������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������GGG�555���������555�999�������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������111�����������������111�nnn���������������������������������������������jjj�[[[�```�����������������UUU�������������������������222�JJJ�����������������JJJ�111���������������������������������������������jjj�[[[�```�����������������UUU���������������������VVV�111�������������������������111�GGG�����������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������jjj�[[[�```�����������������UUU�����������������������������������������������������������������������������������������������������iii�[[[�___�UUU�XXX�XXX�XXX�XXX�XXX�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�YYY�UUU�\\\�fb� 5   b� �������� � ���� � �     X O R   J u n c t i o n 1   X O R   J u n c t i o n [ I D E F 3   p r o c e s s   s c h e m a t i c   s y m b o l s . c d l ] �� ������ pb�       Y@       Y@               ��@      ̐@    �7� J          �?     I@�Y� J          �?      I@ ij�         @�     Y@�����x�      Y@ j��  ���� ���� � �          �v� ����� ݠ ��������p�� �� C   *   W      @�� C   *    X   `U}I@         �-� J          �?     I@�T� B           �?   XU__@    �z� J          �?      @��� J          �?   `U}9@ i�� ��� @   ~         @      @      @   `U�G@     q�      �        ��% % %                   r>�                                             so�     @@   @@   @@   @@ �       �B      �v�      ��� ��� J                ��� J                ��� �֡ J            Y@��� J                �=� �� J                �5� J             Y@�~� �X� J            Y@�v� J             Y@                {��                           ���       |�                                       %�� ����K�  ��     ��               �*�             �����K�    X O R   j u n c t i o n 9�� ������    X O R   J u n c t i o n         ���     ���        <�� ������  =ݣ ����ݣ                       �?      �?                ?� �����  C � ��������                              �?        Z� ��������E� ����E�    fQ� ;   Q� ����Z� ߩ ����<� ǩ ��������k� ���������            ٥ ����� p�� ��� K	            S     Y@�� K	            S      Y@         �� J          �?     I@�<� J          �?      I@    �b� J          �?     I@��� J          �?      I@ i�� ��� A   ~                Y@              Y@ j٥  ���� ���� � �          ��� ����e� (� ��������p� �(� K            S     Y@�R� K            S      Y@         �}� J          �?     I@��� J          �?      I@    �Ŧ J          �?     I@�� J          �?      I@ i� �� @   ~   t�q��@@�qǡ�P@   @U�0@   ���T@     qX�     �        ��% % %                   r��                                           X s�  ��� B    �������?  �A�ϧ B    �������?  �A   @@   @@ �       �B      ���                       {4�                           �4�       |e�                                       %s� ������  �|�     ���               ���             �������     9ݨ ����ݨ             �Ш     �ݨ        <� �����  =(� ����(�                       �?      �?                ?6� ����6�  Ck� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         uǩ   ��    ��                                   m<�      n2� �� k                �*� k                nt� �N� j                �l� j             Y@n�� ��� j            Y@��� j             Y@n�� �Ҫ j            Y@�� j                n<� �� b                  �4� b                  &Q� ��������2       fE� ;   E� ��������Ӯ ����0� �� ��������_� ���������            ۬ ����Y� p�� �˫ G    333333�?     .@��� O	            S      Y@         �� N                �B� N          �?      I@    �d� J                ��� J          �?      I@ i�� ��� @   ~                .@              Y@ j۬  ���� ���� � �          �                     {(�                           �(�       |Y�                                        %g� ������  �p�     ���               ���             �������     9ѭ ����ѭ             �ĭ     �ѭ        <߭ ����߭  =� �����                       �?      �?                ?*� ����*�  C_� ��������                              �?        t��          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                   m0�      n&� � � k                �� k                nh� �B� j                �`� j             Y@n�� ��� j            .@��� j             Y@n� �Ư j            .@�� j                n0� �	� b                  �(� b                  &E� ��������2       V� ��������       �b�   �׺ l
  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  	�IDATx�]g�K���3���E����ADP1��@`�1bΊa�9��&��O�?#��30�j_U���[��{�޺��{�3����	�� ���G��#�sLJJ���ϟ����6g����у��\%7��ٳ瞔��%K���c:�ȧ�/&5m��]L'�F9��Ǐ�322.�.�.r��B�ҩ��I�z���c:fffRZZ�?�HL'�F9�@�KJk׮U������K��N�T<X�D,iW;-"P�`Y��]�@ŃeID��v��"�%K��N�T<X�D,iW;-"P�`Y��]�@ŃeID��v��"�%K��N�T<X�D,iW;-"P�`Y��]�@ŃeID��v��"�%K��N�T<X�D,iW;-"P�`Y��]�@ŃeID��v��"�%K��N�T<X�D,iW;I\�z���h�="u�/_>*_��.���^�zEo߾5��t��T�pac<QN�����4m�4#�y��={�P�*U�ub|������Kϟ?7�b͚5J�g�'j���A۶m�bŊF,�}�F���3��	�`� Z�n� ��S"ȟ??M�4�������ԩS�:��޽K;w�46+X�`��26N��S" ^-Z�����[�[�p!�2wZ�d7����3g�h��#GR�r�L��;' ʘJ���?�Y�v������G7o�4V�_�>ś	�x��pRe˖��Ç[!ڱcݿ�Z'(���KZ�b��Z�ܹi��锜�$������ݻ7լY�WG����Ms��5�Nf��+/^��޿��}��ի��A�\�h�ԩJ�o��ڵkt��c��p���dx2d�)��Y �z��!M��K�Zxt��~����">�W`p�sZ  O�J�2r����}]�p����I]�nݺQ�F�La��΋�H�"4n�8+����[�nY�D��NOO��u�?3f̿�.;���ܹ35i�������#��0�ہ��zZ�hQS�I�" �'O&���Ν;�yS�'NM��*�7�FU�V��Z�Y�j��_g�޽�E��Ba��!4���A�Q�ʕ�<�o:�	�G�A*T�5u������m=v�]�|Y!���6Y�:u�O�>���~�D 6�5kF�:u���?L;�0�8{�l��"�04����@^m+|<x@۶ms�{�n�T�����g�6�s�����H6[�nݸq�V�6�c�J�*�СCm��"����q/7��ϟ	@X6f2�M��w�V����N�v�����bъ�[ �ڵkǴ�x��C���������2e�D�,!.�����^1q+�dދ dv�Ё�7o�+���9���H����
*�Mn�;���nڴ)���/_hٲe��|��� +�222��ݡC���ի٪�K%�E���CڰaCT|a.!2�UCG+{-�(�5kVԄbna�֭�R���Z�+W�D�J������ɓ'1�u���"x��q	HB�5j���BN�p6^�����󭻇�Tlƌֹ��g���ӧ�5��^��̙3V�ڵkG-[��Z�j�-,X��:����ʹ+y'lI���c7�	~!���?0v8#A���V�\IϞ=3r����1�-�;6R���¶�H��!�W"�J�]�v�7M-cH�q���vHP��[�
ccވ �;0e6���)S��"&�L��{��5���{#�-[�X�R �Hݺu�dU�V���Ҍqp����o���GM�?<��� b�m�R��5�p��Dj[�!�@�ʛC����ɓ'	�|2�Ep��a�t钑,&�ر�1�5ЦMjժUV�R��L;�bN� if�W�d�$��P�v�ĉ�,$�?��7�:�sZ�Wh�5<x�`��hO��a���}0gEp�ܹp>	x���X������&����kdj�h~'E��ӧp���%���Em�n%x9z�hЩ>�0����S#�]�v���� cy��%K�XoIٽ֟��n߾M۷o7bV�X1=z�1m �
�ȯ_���˗G{ڄ���K`�̙�1�Q�FQ�%�3��{iذa��!;���׭u9��S�޽{F<4h�1h�c )tSRR����.�S"@�j�a���4���A~lJ	JZ�dڮ.U7O�!��\�9�qRSSc^��ӟ-��;�Kog���V^+����qa���[�Y�V^+����qa���[�Y�V^+����qa���[�Y�V^+����qa���[�Y�V^+����qa���[�Y�V^+����qa���[�Y�V^+����qa���[�Y�V^+������ :�#8C*x����<�|ikG ��)dʗ?	��ݻw	%g:�����89[��9�y!�]"��y\zz�����V�D�o�~�6<fI    IEND�B`�   g2�     .� ����;� 4   C a l l   a n d   C o n t i n u e   R e f e r e n t           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�WWW�~~~�}}}�yyy�yyy���������������������������������������������������������������������������������������������������������ccc�]]]�UUU�����������������UUU�����������������������������������������������������������������������������������������������������UUU�YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�{{{�����������������jjj���������������������������������������������������������������������������������������������������������YYY�UUU�����������������^^^�����������������������������������������������������������������������������������������������������xxx�YYY�VVV�{{{�{{{�{{{�{{{���������������������������������������������������������������������������������������������������������UUU�WWW�{{{�����������������������������������������������������������������������������������������������������������������������������WWW�{{{�����������������������������������������������������������������������������������������������������������������������������WWW�{{{�����������������������������������������������������������������������������������������������������������������������������WWW�WWW�����������������������������������������������������������������������������������������������������������������������������WWW�```�hhh�iii�iii�iii�iii�iii�jjj�jjj�jjj�jjj�jjj�jjj�jjj�kkk�kkk�kkk�kkk�kkk�kkk�lll�lll�lll�lll�lll�mmm�mmm�mmm�mmm�mmm�ggg�aaa�[[[�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f
� 5   
� ��������� ����� 7 �    C a l l   a n d   C o n t i n u e   R e f e r e n t 9   C a l l   a n d   C o n t i n u e   R e f e r e n t [ I D E F 3   r e f e r e n t s   a n d   n o t e s . c d l ] �� ������ p��  ������x@ p�'�Y�o@          �q��G�@      ڢ@    �{� J          �?������h@��� J          �?p�'�Y�_@ i��       ��ư�������x@        p�'�Y�o@ j��  ���� ���� � �          ��� ������ � ��������p�� �(� C    L    P�����t@�J� C        V�oY�g@         �q� J       ������x@��� J                    ��� J       P�����t@��� J                 i�� ��� @   ~         $@    R�o@      $@   ���W@     q@�     �      
  ��% % %                   rq�                                            R e f e r e n t   T y p e /   L a b e l s��       A    A    A    A �       �B      ���      �� ��� J                �� J                �W� �1� J                �O� J       p�'�Y�o@��� �r� J       ������x@��� J                ��� ��� J       ������x@��� J       p�'�Y�o@   }`� ��� C       �Q� @P@�� G        V�oY�g@�4� B   L    �Q� @P@�O� B   M    V�oY�g@           d?� ��� B   L        
   	      C o n t r o l s . x 1       Y               �7� B   L     333333�?         C o n t r o l s . x 1  333333�?  Y                       {r�                           �r�       |��                                       %�� ���� �  ���     ���               ���             ����� �    c a l l   a n d   c o n t i n u e   r e f e r e n t 9�� ������ 4   C a l l   a n d   C o n t i n u e   R e f e r e n t         �v�     ���        <�� ������  =�� ������                       �?      �?                ?�� ������  C� ��������                              �?        � ���������� ������    f8� ;   8� ����A� �� ����#� �� ��������N� ��������8            �� ����H� p~� ��� O	            S������x@��� O	            Sp�'�Y�o@         �
� N          �?������h@�-� N          �?p�'�Y�_@    �S� J          �?������h@�u� J          �?p�'�Y�_@ i�� ��� @   ~   {�b#�ư�������x@        p�'�Y�o@ j��  ���� ���� � �          �                     {�                           ��       |H�                                        %V� ������  �_�     �s�               ���             �������     9�� ������             ���     ���        <�� ������  =� �����                       �?      �?                ?� �����  CN� ��������                              �?        tr�          ��U U U          �?u��   ��  ��� � �         u��   ��    ��                                    m#�      n� ��� k                �� k                n[� �5� j    � ��D=fiI�M��=�S� j       p�'�Y�o@n�� �w� j       ������x@��� j       p�'�Y�o@n�� ��� j       ������x@��� j                n#� ��� b                  �� b                  &8� ��������2       f� ;   � ����� �� ������ �� ��������&� ��������9            �� ������ pn� ��� G       ������x@��� K	         �{��S�?S�Q� @P@         �� N                �%� N       p�'�Y�o@    �G� J                �e� J       �Q� @P@ i�� ��� A   ~   {�b#�ư�������x@        �Q� @P@ j��  ���� ���� � �          ��� ���� � 	� ��������p�� �	� K            S������x@�3� K            S�Q� @P@         �^� J          �?������h@��� J          �?�Q� @@@    ��� J          �?������h@��� J          �?�Q� @@@ i�� ��� @   ~   ��8�I�a@8��8[p@�zDa��&@�Q�U�J@     q9�     �      
  ��% % %                   rj�                                           L o c a t o r s��      A    A    A    A �       �B      ���                       {��                           ���       | �                                        %.� ����i�  �7�     �K�               �`�             �����i�     9�� ������             ���     ���        <�� ������  =�� ������                       �?      �?                ?�� ������  C&� ��������                              �?        tJ�          ��U U U          �?uh�   ��  ��� � �         u��   ��    ��                                    m��      n�� ��� k                ��� k                n3� �� j    � ��D=fiI�M��=�+� j       �Q� @P@nu� �O� j       ������x@�m� j       �Q� @P@n�� ��� j       ������x@��� j                n�� ��� b                  ��� b                  &� ��������2       f�� ;   �� ��������{� ������ c� ��������� ��������5            �� ����� p7� ��� G   L    �Q� @P@��� G        V�oY�g@         ��� N                ��� N                    �� J                �.� J                 iN� �L� @   ~   ���ư��Q� @P@        V�oY�g@ j��  ���� ���� � �          �                     {��                           ���       |�                                        %� ����J�  ��     �,�               �A�             �����J�     9y� ����y�             �l�     �y�        <�� ������  =�� ������                       �?      �?                ?�� ������  C� ��������                              �?        t+�          ��U U U          �?uI�   ��  ��� � �         uc�   ��    ��                                   m��      n�� ��� k                ��� k                n� ��� j                �� j       V�oY�g@nR� �,� j       �Q� @P@�J� j       V�oY�g@n�� �n� j       �Q� @P@��� j                n�� ��� b                  ��� b                  &�� ��������2       �� ��������       �
�   �.�   �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�KH\Y��:�Zc4$>��J�E&>����F	�WA]h@	�
YJp!���5���"b��&�r�M��czn��gp1]���4�m��~�ϩ{{!� � � � � � � � � � � � � � � � � � � � � � � �N���e+--����|��aaa���H�����z{{�����X���=�'M�pyR�{��(�Y!!!����r:��U�tww��k��QGGG���P�B !��`�� \-����D�j�F�8%X'B W�4B��)�:A�Z�-N	։��"�hqJ�N�@�i�@�S�u"�p�H#Z��!��E!��`�� \-����D�j�F�8%X'B W�4B��)�:A�Z�-N	։��"�hqJ�N�@�i�@�S�u"�p�H#Z��!��E!��`�� \-����D�j�F�8%X'B W�4B��)�:A�Z�-N	։��"�hqJ�N�@�i�@�S�u"�p�H#Z��!��E!��`�� \-����D�j�F�8%X'B W�4B��)�:A�Z�-N	�iݿ�g�_��f��\�M���K�.]��� �iB��������o��6�{�=z���lYEDDx�j(z���������Ϫ��������	 ������������!G�� ��x��8b�@u���hkk��){y��CP[[K/_��8���Y*((𸮷
�}��՝�.�	233CGGG���N�/_6J����^=RSSͽ�ׯ_Ӈ�o�edd��奥%��ߧ��y
		���$ZYY!~�k�(--��^ț7oȾ�F��666(>>�����|.���R�����cypp@]]]H��崺�J7nܠ��z��)555��o߾5Ntwwӳg�h{{�ZZZ���딗�G555���L���t��]z��	������2qh�������|�<��>���	s�vtt�-Q������s���������Y�f������ }��޽{GEEE�Ъ�*��R{{��ZWWG<0Z�߿���B�����������h����B0::J����ƿ����U�Ν;�4��g8���c����+W��0�6pr|��^�xAeee�e6;!!�����s�n4���BF��{�����U�mmm潼:�w����v�\�w��'5Y�� ���M�{}}�<�9��ͥ��IӴ����U����7oo�a���3!���"pm.=Y�W�L�X��������_	��ી��aJII���b��ߺu�rrr�����+���W�������Ç����s�Ϗ��8�}�6ݻw�hqP]]mD�⨬�4�O���>����t�L�v:�����*�p��������3ܽ�s����G�$�����Mc6_Y����cxx�q �%�����uvv��s=��n�N����=xo����wHLL���O�T����t0�9���i�v`w�w�� �Fv�cY������ﮝ��^,.�h��R����B4@ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @�+�!����    IEND�B`�   gI"     E" ����R" ,   C a l l   a n d   W a i t   R e f e r e n t           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�]]]�������������������������������������������������������������������������������������������������������������������������lll�]]]�]]]�������������������������������������������������������������������������������������������������������������������������mmm�]]]�]]]�������������������������������������������������������������������������������������������������������������������������nnn�]]]�[[[�������������������������������������������������������������������������������������������������������������������������hhh�]]]�UUU�ddd�ddd�ddd�aaa�___�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�kkk�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�jjj�aaa�```�ddd�ddd�ddd�UUU�YYY���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX���������������������qqq���������������������������������������������������������������������������������xxx���������������������XXX�vvv�����������������nnn���������������������������������������������������������������������������������ppp���������������������XXX�UUU�]]]�]]]�]]]�XXX�ccc�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ggg�ccc�[[[�]]]�]]]�]]]�UUU�WWW���������������������������������������������������������������������������������������������������������������������������������XXX���������������������������������������������������������������������������������������������������������������������������������XXX���������������������������������������������������������������������������������������������������������������������������������XXX���������������������������������������������������������������������������������������������������������������������������������XXX�UUU�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�WWW�UUU�YYY�[[[�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f! 5   ! ��������O ����O � �    C a l l   a n d   W a i t   R e f e r e n t 5   C a l l   a n d   W a i t   R e f e r e n t [ I D E F 3   r e f e r e n t s   a n d   n o t e s . c d l ] "� ����0� p��  ������x@ p�'�Y�o@          gffff��@ wwwwwa�@    ��� J          �?������h@��� J          �?p�'�Y�_@ i��    �=#K��������x@T����1��p�'�Y�o@ j"�  ���� ���� � �          � ����� ^  ��������p&  �n� C    L       �p׫��p@��� C        V�oY�g@         ��� J          �?������h@��� J                    ��� J          �?�p׫��`@�  J                 i<  �:  @   ~         $@    R�o@      $@   ���W@     q�      �      
  ��% % %                   r�                                             R e f e r e n t   T y p e /   L a b e l s       A    A    A    A �       �B      �      �d �> J                �\ J                �� � J                �� J       p�'�Y�o@�� �� J       ������x@�� J                �' � J       ������x@� J       p�'�Y�o@   }� �E C       �Q� @P@�g G        V�oY�g@�� B   L    �Q� @P@�� B   M    V�oY�g@           d� � B   L        
   	      C o n t r o l s . x 1       Y               �� B   L     333333�?         C o n t r o l s . x 1  333333�?  Y                       {�                           ��       |�                                       %� ����f  �     �               �1             �����f    c a l l   a n d   w a i t   r e f e r e n t 9� ����� ,   C a l l   a n d   W a i t   R e f e r e n t         ��     ��        <� �����  = ����                       �?      �?                ? ����  CO ��������                              �?         �������� ����    fv
 ;   v
 ����
  	 ����a
 � ��������� ���������             ����� p� �� O	            S������x@� O	            Sp�'�Y�o@         �H N          �?������h@�k N          �?p�'�Y�_@    �� J          �?������h@�� J          �?p�'�Y�_@ i� �� @   ~           ������x@        p�'�Y�o@ j  ���� ���� � �          �                     {U                           �U       |�                                        %� �����  ��     ��               ��             ������     9� �����             ��     ��        < ����  =I ����I                       �?      �?                ?W ����W  C� ��������                              �?        t�          ��U U U          �?u�   ��  ��� � �         u�   ��    ��                                    ma
      nS	 �-	 k                �K	 k                n�	 �s	 j    � ��D=fiI�M��=��	 j       p�'�Y�o@n�	 ��	 j       ������x@��	 j       p�'�Y�o@n
 ��	 j       ������x@�
 j                na
 �:
 b                  �Y
 b                  &v
 ��������2       fN ;   N ����W � ����9 � ��������d ���������            � ���� p� ��
 G       ������x@� K	         �{��S�?S�Q� @P@         �D N                �c N       p�'�Y�o@    �� J                �� J       �Q� @P@ i� �� A   ~           ������x@        �Q� @P@ j�  ���� ���� � �          �� ����^ G ��������p �G K            S������x@�q K            S�Q� @P@         �� J          �?������h@�� J          �?�Q� @@@    �� J          �?������h@� J          �?�Q� @@@ i% �# @   ~   ��8�I�a@8��8[p@�zDa��&@�Q�U�J@     qw     �      
  ��% % %                   r�                                           L o c a t o r s�      A    A    A    A �       �B      ��                       {-                           �-       |^                                        %l �����  �u     ��               ��             ������     9� �����             ��     ��        <� �����  =! ����!                       �?      �?                ?/ ����/  Cd ��������                              �?        t�          ��U U U          �?u�   ��  ��� � �         u�   ��    ��                                    m9      n+ � k                �# k                nq �K j    � ��D=fiI�M��=�i j       �Q� @P@n� �� j       ������x@�� j       �Q� @P@n� �� j       ������x@�� j                n9 � b                  �1 b                  &N ��������2       f+ ;   + ����4 � ���� � ��������E ��������0            � ����? pu �� G   L    �Q� @P@�� G        V�oY�g@         � N                �, N                    �N J                �l J                 i� �� @   ~           �Q� @P@        V�oY�g@ j�  ���� ���� � �          �                     {                           �       |?                                        %M �����  �V     �j               �             ������     9� �����             ��     ��        <� �����  = ����                       �?      �?                ? ����  CE ��������                              �?        ti          ��U U U          �?u�   ��  ��� � �         u�   ��    ��                                   m      n �� k                � k                nN �( j                �F j       V�oY�g@n� �j j       �Q� @P@�� j       V�oY�g@n� �� j       �Q� @P@�� j                n �� b                  � b                  &+ ��������2       f ;    ��������� ����� z �������� ��������1            � ���� pN �� G       �Q� @P@�� G       V�oY�g@         �� N       ������x@� N                    �' J       �Q� @P@�E J                 ie �c @   ~           �Q� @P@        V�oY�g@ j�  ���� ���� � �          �                     {�                           ��       |                                        %& ����a  �/     �C               �X             �����a     9� �����             ��     ��        <� �����  =� �����                       �?      �?                ?� �����  C ��������                              �?        tB          ��U U U          �?u`   ��  ��� � �         uz   ��    ��                                   m�      n� �� k                �� k                n' � j                � j       V�oY�g@ni �C j       �Q� @P@�a j       V�oY�g@n� �� j       �Q� @P@�� j                n� �� b                  �� b                  & ��������2        ��������       �!   �E"   �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  �IDATx�_H�Y���X�i�n%�F�2����+1��<"Q>H(؃�(�>mAD=���(F� ��&X+�b��R0m���߹����&P�㙙�����3���w����� � � � � � � � � � � � � � � � � � � � � � � �p���D�\�^����}���i�v8�]��l	X<�-�	�'�h��kjj��K��766�*++�����v�x<���t�h�7�����|L�:::�����9�����m��{bߕ������v��+@4����������>��}vv����(h�N�3�	���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S���&��=L�]!��`��S�oH;����Z���hxx����3�-//�Ǐ)�:qL>�֗&�������?h�O�<I�N������Ō�@�Lt��ՠ������u�i}������>��aNkkk�[ߕ�#Lx���Q��6� ��{�0��kY���қ7o"L��y�!k���q���=*�?��O�Il�A�f���SӧO��ݻw���L999d=�p_�|��oߚ=�k׮�v�H����v�iss�>�LQQQ4::J)))t��9��i=g�X111�/�)�خ;R}}=eff���$ݸq�=zDCCC���H�ϟ7���ѝ;w����\.���Z[[���8l�۷oә3glc>�����ijj��_�NϞ=;6!�8�L���EUUUTSSc���^��K�<yB�nݢ�`bb�.^�H������m����2:}�4y<�]Ԧ�&Ö���<��|�Ҍ��8��5���߿��� ����<��Я^�2��͛7w��+W��;�G����w�1÷o��:P̝m���ܐ6 �ٰ	�N'������+���:��Ǜ)`o;w��MMߞ�JHH������x���@1y��#�G��r��w1�|>���_�6��N��Φ��N���ʊ��:-���̧�;&�p�����y$�����.ݑ�n��/))������޽KuuuTXXH[[[t��}3:�����JKKͰ�>~544����Wqq1�x�´�ch�������ᨨ�h����5�>E䡜�Ξ=k�W$^���S_�~%RSS�'(������G1�������3��;���C�����=xn4�'%%�v�Q��N!�Kȯ	B����aUrO10��pW��i����hZ]]�σ���P�Q���R�1b�o��ҟ�d	G�����a=
���2T                                         ����+k��� t�    IEND�B`�   gTM     PM ��������   N o t e           �?�   !   !                                                                                                                                       ����]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�]]]�����]]]�������������������������������������������������������������������������������������������������������������������������jjj�]]]�ZZZ�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�yyy�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�xxx�yyy�xxx�xxx�yyy�yyy�xxx�xxx�www�aaa�[[[�����������������������������������������������������������������������������������������������������������������������������UUU�[[[�����������������������������������������������������������������������������������������������������������������������������___�[[[���������}}}�����������������������������������������������������������������������������������������������������������������___�[[[�������������yyy�������������������������������������������������������������������������������������������������������������___�[[[�mmm�}}}�}}}�}}}�}}}�|||�|||�}}}�|||�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�}}}�UUU�[[[�����������������������������������������������������������������������������������������������������������������������������^^^�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�����������������������������������������������������������������������������������������������������������������������������```�\\\�\\\�|||���������������������������������������������������������������������������������������������������������������������```�\\\�\\\�����|||�����������������������������������������������������������������������������������������������������������������```�\\\�]]]���������|||�������������������������������������������������������������������������������������������������������������```�\\\�]]]�������������}}}���������������������������������������������������������������������������������������������������������```�\\\�]]]�����������������}}}�����������������������������������������������������������������������������������������������������```�\\\�]]]���������������������ooo�}}}�~~~����������������������������������������������������������������|||�UUU�\\\�]]]��������������������������������������������������������������������������������������������������������������������������]]]�]]]�����������������������������������������������������������������������������������������������������������������������������]]]�]]]�jjj�lll�mmm�nnn�ooo�ppp�rrr�sss�uuu�vvv�www�www�xxx�yyy�{{{�|||�}}}�~~~��������������������������������������������������]]]�f~D 5   ~D �������� 8 ���� 8 M �    N o t e #   N o t e [ I D E F 3   r e f e r e n t s   a n d   n o t e s . c d l ] �4 �����4 p�4        t@ ���T�Jp@          �i����@ �NTx!�@    �e4 H          �?      d@��4 H          �?���T�J`@ i�4                  t@        ���T�Jp@            ��6 ����
7 6 ��������p�5 �5 H          �?         S      t@�35 C        XUU@�j@         �^5 H          �?      d@�|5 J       ���T�Jp@    ��5 H          �?      d@��5 J       XUU@�j@ i�5 ��5 @   ~         4@      4@      4@   ��*O@     q16      �      
  ��% % %                   rb6                                              s�6      �A   �A   �A   �A �       �B      ��6                       {�6                           ��6       |
7                                       %7 ����[7  �!7     �57               �J7             �����[7    n o t e 9�7 �����7    N o t e         ��7     ��7        <�7 �����7  =�7 �����7                       �?      �?                ?�7 �����7  C 8 ��������                              �?        vD ��������aD ����aD    f�= ;   �= �����= �; ����r= �; ��������J; ��������K            �9 ����D: p�9 ��8 O	            S      t@��8 O	            S���T�Jp@         �9 N          �?      d@�<9 N          �?���T�J`@    �b9 J          �?      d@��9 J          �?���T�J`@ i�9 ��9 @   ~                 t@        ���T�Jp@            �                     {:                           �:       |D:                                        %R: �����:  �[:     �o:               ��:             ������:     9�: �����:             ��:     ��:        <�: �����:  =; ����;                       �?      �?                ?; ����;  CJ; ��������                              �?        tn;          ��U U U          �?u�;   ��  ��� � �         u�;   ��    ��                                   mr=      n< ��; k                �	< k                n`< �-< j                �X< b         @P@ | XUU��uh@n�< ��< b        @P@ |      @P@��< j       ���T�Jp@n�< ��< j             t@��< j       ���T�Jp@n.= �= j             t@�&= j                nr= �K= b                  �j= b                  &�= ��������2       faD ;   aD ���������B ����LD �B ��������{B ��������L            ? ����? p�> �
> K	            S      t@�+> C   *    X   ��*H@         �W> N          �?      d@�v> N                    ��> J          �?      d@��> J                 i�> ��> A   ~                 t@           ��*H@ j?  ���� ���� � �          �A ����uA ^@ ��������p&@ �^? K            S      t@��? K            S   ��*H@         ��? J          �?      d@��? J          �?   ��*8@    ��? J          �?      d@�@ J          �?   ��*8@ i<@ �:@ @   ~         4@����̥a@      @   ���F@     q�@     �      
  ��% % %                   r�@                                            N o t e   I D s�@     �A   �A   @@   @@ �       �B      �A                       {DA                           �DA       |uA                                        %�A �����A  ��A     ��A               ��A             ������A     9�A �����A             ��A     ��A        <�A �����A  =8B ����8B                       �?      �?                ?FB ����FB  C{B ��������                              �?        t�B          ��U U U          �?u�B   ��  ��� � �         u�B   ��    ��                                   mLD      nBC �C k                �:C k                n�C �^C j                �|C j          ��*H@n�C ��C j             t@��C j          ��*H@nD ��C j             t@� D j                nLD �%D b                  �DD b                  &aD ��������2       rD ��������       �~D   �PM �  �PNG

   IHDR   �   �   ��P   sRGB ���   DeXIfMM *    �i            �       �       ��       �    �H�  3IDATx�klL[�׌I+�{����x�z4�􁆐ho�����F�7��M<>�E$�	M�$hBI�H)q[7��h�Ѫ>�Y���i;��5��۳�?pz�^{�������� � � � � � � � � � � � �p��3�n��~�qj/_�\�Z�hQv�n�
z���y#K�ϟ?�$��f��	&4�ڵ��
��[?�cǎ5��������C����uHE��'T����@ֳ�t��Ƞ��xs�;?n�8�ׯ�9�?���������.���O�NO�<�O�>�ܽ{w�ի�5��Ů��	�%����i˖-f�͛7��ի�q}}�9�w�^�7o^�O����Y�f��ݻiΜ9A�����W:r����������	���Z��������7��ٳ�s���m;s���ֶ&�������jjj
�9@�>}�����i�ȑ���J׮]�{�;�=zD�nݢ�Ǐ�ݹs�={�q��H�5k�З/_���0�`,����7033�|+++M_�L��\�СC���{��̒��N���'��E��C�����Q��8q�F�A;v����P�1]$��a�(++�Ξ=K߾}koϞ=��\��+Wҳg�hݺu���)S���cƌ��3g��ɓ��ÇF��'��Çiڴit��z��A��%'hŊ��z���L�}E0������Z �����7o���߰a�۷�<�oܸA,0��N�J�����g�%x����KÇ����cG�/����FS1a-��2�,

h�ܹ��ׯ_��I�&�����4_�b�n�^�2ח-[f_b�xa���[����Xn���t��U:��=:������>�[I�����:�Wִ|���y����RRR::����$0` �汅�6�?~L����ӧ�àA��};�[�5�U޼yC3f�0�|�y�It����өS����ZpI�C�]���\�bF��3x���t��%JJJ2S�ɓ'�~?��2��m\rr��f����[��x�� ��>¿����˗f��k���8�����/^�0�Ǟ={��
�c�80��������KK�.�s����b.����i�����W�,7�=z�������-UWWS~~>ݾ}��ILL�M�6�c�?>|�@�V�2�޾}k��n�[EEm۶�<�X�ŋ���}��?�%�Z�d��ִ�[g�*��[ȡC��5���󾝯�4���� �$�޽3{������q������L���,�^�w����o<ô>���%`$��m{+��~<F�?	��K���ϟ��y�[��/���XSq��&��~�[���&�Z�D�B������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*������j*��m��I��_�(�D�n��[XZZZ���W�&+$""�.**����c�ݻw��"vj:�5DPSψ��!"~*�l	8�����$ZH�J��ӧOc�(F꼀6���^RR�WS�� "�9::�]	 ���*���@K�v)Dplmþ�$�a�tdǰ%���oX7-� "���q��@��8�G$D��Q"� "8��Ao�C@��ls��@�Ժ��	 B�|q��$���w���T	Z�P�����{�:�����v���е��n�"DȺ˞����ּ͍�ڜ�����ѣG�QYY���x��2qMMM���?��e��K���(HHHh�x���QÂ � � � � � � � � 8��?'����    IEND�B`�   	iM ����iM     �����M �����M   ��       ��� � � ��          �      T a h o m a ����    ��M     ��M     -�M �������� � Q                  �}N                               	   
                                                          S e c t i o n   1 ��N                     ��N                     ��N                     ��N                     ��N                     �O                     �,O                     �EO                     �^O                     �wO                     ��O                     ��O                     ��O                     ��O                     ��O                     �P                     �&P                     �?P                     �XP                     �qP                     ��P                     ��P                     ��P                     ��P                     ��P                     �Q                     � Q                     